
`timescale 1ns / 1ps

module tb_N8_restoring_divider;

    // Parameters
    
    parameter N = 8;
    
     
    // Inputs
    
    reg   clk;
    
    reg   rst;
    
    reg   start;
    
    reg  [7:0] X;
    
    reg  [7:0] Y;
    
    
    // Outputs
    
    wire  [7:0] quot;
    
    wire  [7:0] rem;
    
    wire   valid;
    
    
    // Instantiate the Unit Under Test (UUT)
    restoring_divider  #( N ) uut (
        
        .clk(clk),
        
        .rst(rst),
        
        .start(start),
        
        .X(X),
        
        .Y(Y),
        
        
        .quot(quot),
        
        .rem(rem),
        
        .valid(valid)
        
    );

    // Clock generation 
    
    
            always begin
                #5 clk = ~clk;
            end
            
    

    
    
            always begin
                #99 rst = 1'b1; 
            end
            
    
    
    initial begin
        // Initialize Inputs
        
        clk = 0;
        
        rst = 0;
        
        start = 0;
        
        X = 0;
        
        Y = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 X = 8'b00100000; Y = 8'b11001001; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 0,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b00111100; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00010001; // Expected: {'quot': 3, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 3,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b01101111; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 4,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10001000; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 5,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b01100101; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 6,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 7,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 8,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 9,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b01110000; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 10,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 11,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00001010; // Expected: {'quot': 4, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 12,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b01111011; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 13,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 14,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 15,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b00101010; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 16,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 17,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b00111100; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 18,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b01001000; // Expected: {'quot': 2, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 19,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b10100011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 20,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 21,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10011011; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 22,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 23,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b01111100; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 24,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00111011; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 25,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b00111010; // Expected: {'quot': 3, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 26,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 27,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 28,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 29,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b01101110; // Expected: {'quot': 1, 'rem': 105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 30,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11100101; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 31,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 32,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 33,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b01011111; // Expected: {'quot': 2, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 34,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b11011000; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 35,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01100000; // Expected: {'quot': 1, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 36,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b00011101; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b00011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 37,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 38,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 39,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 40,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 41,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01111111; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 42,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00101101; // Expected: {'quot': 3, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 43,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 44,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b01010000; // Expected: {'quot': 1, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 45,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00001010; // Expected: {'quot': 24, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 46,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 24, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10111011; // Expected: {'quot': 1, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 47,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10100001; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 48,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 49,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 50,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 51,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10000110; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 52,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01000110; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 53,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00001101; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 54,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 55,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00101100; // Expected: {'quot': 2, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 56,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00100001; // Expected: {'quot': 2, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 57,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00001100; // Expected: {'quot': 3, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 58,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 59,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 60,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b00010000; // Expected: {'quot': 15, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 61,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b10011110; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 62,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 63,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01000100; // Expected: {'quot': 2, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 64,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b01000010; // Expected: {'quot': 1, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 65,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01001100; // Expected: {'quot': 1, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 66,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 67,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b00111101; // Expected: {'quot': 3, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 68,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01011111; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 69,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b01100001; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 70,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01100011; // Expected: {'quot': 1, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 71,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 72,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b11001100; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 73,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b00101111; // Expected: {'quot': 3, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 74,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10001111; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 75,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 76,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 77,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b01011001; // Expected: {'quot': 2, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 78,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b10100100; // Expected: {'quot': 1, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b10100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 79,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b01011101; // Expected: {'quot': 2, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 80,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b00000110; // Expected: {'quot': 13, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 81,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 82,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 83,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b01111110; // Expected: {'quot': 1, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 84,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01100101; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 85,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b00111110; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 86,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 87,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b01111100; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 88,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b00001100; // Expected: {'quot': 12, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 89,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b00010101; // Expected: {'quot': 8, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 90,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b01101011; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 91,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b10010010; // Expected: {'quot': 0, 'rem': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 92,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 93,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 94,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b10011000; // Expected: {'quot': 1, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 95,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 96,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b01100111; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 97,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 98,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10001011; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 99,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01000001; // Expected: {'quot': 3, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 100,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b01010110; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 101,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 102,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b10000010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 103,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 104,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b00101010; // Expected: {'quot': 3, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 105,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b10110111; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 106,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 107,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 197}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 108,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b00001101; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 109,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b00011101; // Expected: {'quot': 4, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b00011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 110,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b00011010; // Expected: {'quot': 6, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 111,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01001100; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 112,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01101011; // Expected: {'quot': 1, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 113,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b10011101; // Expected: {'quot': 0, 'rem': 137}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 114,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00001000; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 115,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 116,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 117,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b10001010; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 118,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b10100010; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 119,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 120,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 121,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 122,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b01001101; // Expected: {'quot': 2, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 123,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 124,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b10001000; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 125,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 126,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b00111011; // Expected: {'quot': 3, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 127,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01100100; // Expected: {'quot': 1, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 128,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b01000010; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 129,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b11001110; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 130,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 131,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b01110011; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 132,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 133,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01110001; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 134,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b00100111; // Expected: {'quot': 5, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 135,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00001110; // Expected: {'quot': 13, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 136,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 137,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 160}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 138,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 196}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 139,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00001100; // Expected: {'quot': 17, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 140,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 141,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 142,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01100111; // Expected: {'quot': 1, 'rem': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 143,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 144,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 145,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b01001100; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 146,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10010110; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 147,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 148,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 149,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01111000; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 150,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b00001110; // Expected: {'quot': 16, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 151,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 16, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00110011; // Expected: {'quot': 3, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 152,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b01000110; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 153,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b00111110; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 154,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10001100; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 155,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b01111101; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b01111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 156,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01000000; // Expected: {'quot': 2, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 157,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 158,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 159,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 160,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 161,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 169}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 162,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b11001000; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 163,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01010101; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 164,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 165,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01001010; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 166,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b01011010; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 167,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b01110010; // Expected: {'quot': 1, 'rem': 111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b01110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 168,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 172}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 169,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 170,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 171,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00010001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 172,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b00010101; // Expected: {'quot': 10, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 173,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01010000; // Expected: {'quot': 2, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 174,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b01011100; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 175,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b11000111; // Expected: {'quot': 1, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 176,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11000100; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 177,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b00101111; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 178,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00101100; // Expected: {'quot': 4, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 179,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b01000100; // Expected: {'quot': 2, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 180,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b11011111; // Expected: {'quot': 1, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 181,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11000101; // Expected: {'quot': 0, 'rem': 169}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 182,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00011111; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 183,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01000010; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 184,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00100100; // Expected: {'quot': 2, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 185,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 186,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10011101; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 187,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 188,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b10011101; // Expected: {'quot': 0, 'rem': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 189,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11010100; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 190,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 191,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 192,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 193,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b11110010; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 194,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b00110001; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 195,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 196,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 197,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b00110010; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 198,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b00010000; // Expected: {'quot': 10, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 199,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b10010111; // Expected: {'quot': 0, 'rem': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 200,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11000101; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 201,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b00011010; // Expected: {'quot': 4, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 202,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10000001; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 203,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01110101; // Expected: {'quot': 2, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 204,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 205,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b01110011; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 206,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 207,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 208,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 209,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 213}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 210,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 200}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 211,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b01011100; // Expected: {'quot': 2, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 212,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b00001111; // Expected: {'quot': 7, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 213,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10111001; // Expected: {'quot': 1, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 214,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01101011; // Expected: {'quot': 1, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 215,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b11100000; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 216,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 217,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 218,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b01111101; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b01111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 219,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 218}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 220,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b10011000; // Expected: {'quot': 0, 'rem': 133}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 221,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10110011; // Expected: {'quot': 1, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 222,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11101011; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 223,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b01111001; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 224,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 225,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 226,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01001011; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 227,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 228,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 229,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b00111000; // Expected: {'quot': 2, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 230,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b01000101; // Expected: {'quot': 1, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 231,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 232,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 233,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b01101110; // Expected: {'quot': 1, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 234,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 235,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01000101; // Expected: {'quot': 2, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 236,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 237,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00101111; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 238,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 239,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b00111111; // Expected: {'quot': 2, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 240,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 241,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 242,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b00001100; // Expected: {'quot': 19, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 243,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 19, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 244,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 245,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 246,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 247,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01000111; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 248,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b01100111; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 249,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10010001; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 250,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b00011011; // Expected: {'quot': 7, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 251,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 252,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b11111100; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 253,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00011110; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 254,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 255,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b10010111; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 256,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 257,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b01001101; // Expected: {'quot': 2, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 258,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 259,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b00000010; // Expected: {'quot': 25, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 260,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 261,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b00101110; // Expected: {'quot': 2, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 262,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b00011111; // Expected: {'quot': 3, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 263,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 264,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00111100; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 265,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b10001001; // Expected: {'quot': 0, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 266,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10111000; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 267,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11110111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 268,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01111001; // Expected: {'quot': 1, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 269,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00001110; // Expected: {'quot': 4, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 270,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10011000; // Expected: {'quot': 1, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 271,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01111110; // Expected: {'quot': 1, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 272,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 273,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10100011; // Expected: {'quot': 0, 'rem': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 274,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b01100100; // Expected: {'quot': 1, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 275,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b00010011; // Expected: {'quot': 5, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 276,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b00000110; // Expected: {'quot': 42, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 277,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 42, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00011011; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 278,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 191}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 279,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 280,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 281,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b00111110; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 282,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 201}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 283,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b10111011; // Expected: {'quot': 0, 'rem': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 284,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b10111011; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 285,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 286,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 287,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 288,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00001110; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 289,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b01010110; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 290,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10101000; // Expected: {'quot': 1, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 291,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 292,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00010110; // Expected: {'quot': 3, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 293,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 294,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00111101; // Expected: {'quot': 3, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 295,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 296,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10111011; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 297,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 298,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 299,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b00010101; // Expected: {'quot': 11, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 300,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10100011; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 301,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 302,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10010100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 303,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b00011111; // Expected: {'quot': 2, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 304,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 305,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 306,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 307,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00011111; // Expected: {'quot': 8, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 308,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 309,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b01001011; // Expected: {'quot': 2, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b01001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 310,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b10011000; // Expected: {'quot': 0, 'rem': 137}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 311,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01011100; // Expected: {'quot': 2, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 312,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 313,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b01100100; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 314,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 315,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b01000000; // Expected: {'quot': 2, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 316,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10011111; // Expected: {'quot': 1, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 317,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10100110; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 318,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00100111; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 319,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b10001001; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 320,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 321,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b00011100; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 322,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 323,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b11000001; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 324,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b00101111; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 325,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01111001; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 326,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01010000; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 327,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01000001; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 328,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b01101111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 329,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 330,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 197}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 331,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00101111; // Expected: {'quot': 2, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 332,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 333,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 234}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 334,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01110001; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 335,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00010011; // Expected: {'quot': 11, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 336,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01000001; // Expected: {'quot': 2, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 337,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b10000101; // Expected: {'quot': 0, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 338,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00011110; // Expected: {'quot': 3, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 339,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 340,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 341,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00000110; // Expected: {'quot': 4, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 342,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b11111101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 343,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 344,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01000100; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 345,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01001111; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 346,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 347,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00010110; // Expected: {'quot': 9, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 348,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 349,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01000000; // Expected: {'quot': 2, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 350,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00010001; // Expected: {'quot': 11, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 351,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b00010011; // Expected: {'quot': 3, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 352,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b01011001; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 353,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 354,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b01000110; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 355,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b01100000; // Expected: {'quot': 1, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 356,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01011001; // Expected: {'quot': 2, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 357,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b00111000; // Expected: {'quot': 3, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 358,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 359,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b01010011; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 360,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00100111; // Expected: {'quot': 5, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 361,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 362,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 363,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00101101; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 364,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10110011; // Expected: {'quot': 1, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 365,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 366,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 367,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b10001100; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 368,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00111111; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 369,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01001000; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 370,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00000010; // Expected: {'quot': 113, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 371,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 113, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b00011011; // Expected: {'quot': 2, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 372,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10010011; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 373,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b01111001; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 374,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 375,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b00100010; // Expected: {'quot': 7, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 376,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b10100101; // Expected: {'quot': 1, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 377,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b00100100; // Expected: {'quot': 5, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 378,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b00011100; // Expected: {'quot': 4, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 379,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 380,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 381,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00011010; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 382,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 383,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b00011100; // Expected: {'quot': 3, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 384,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00010110; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 385,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 386,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 387,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b00100010; // Expected: {'quot': 2, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 388,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10011110; // Expected: {'quot': 1, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 389,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00000110; // Expected: {'quot': 34, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 390,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 34, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 391,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b01000010; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 392,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 191}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 393,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00001000; // Expected: {'quot': 5, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 394,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10000111; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 395,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b00110111; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b00110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 396,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 397,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b00011001; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b00011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 398,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 399,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 400,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01010100; // Expected: {'quot': 2, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 401,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 127}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 402,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 403,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00100100; // Expected: {'quot': 5, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 404,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 405,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b00100101; // Expected: {'quot': 6, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 406,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01111100; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 407,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00100111; // Expected: {'quot': 4, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 408,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b01100111; // Expected: {'quot': 1, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 409,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 410,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11010010; // Expected: {'quot': 1, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 411,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 412,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b00100011; // Expected: {'quot': 3, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 413,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b10111100; // Expected: {'quot': 0, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b10111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 414,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b00110010; // Expected: {'quot': 4, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 415,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00110001; // Expected: {'quot': 2, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 416,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10110100; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 417,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b00010010; // Expected: {'quot': 2, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b00010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 418,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 419,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01010101; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 420,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00101000; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 421,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 422,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b00011010; // Expected: {'quot': 4, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 423,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10100101; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 424,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b00100011; // Expected: {'quot': 4, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 425,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b11000001; // Expected: {'quot': 1, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 426,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b10010100; // Expected: {'quot': 1, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 427,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 428,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01111111; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 429,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 137}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 430,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01011101; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 431,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b10010101; // Expected: {'quot': 0, 'rem': 134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b10010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 432,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b01000100; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 433,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 434,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10010011; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 435,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 109}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 436,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11010011; // Expected: {'quot': 0, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 437,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 438,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b01001100; // Expected: {'quot': 2, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 439,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00110001; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 440,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10000111; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 441,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b00111110; // Expected: {'quot': 3, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 442,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 443,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01010000; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 444,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 445,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00001110; // Expected: {'quot': 6, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 446,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 447,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b01001000; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 448,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 449,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b10011111; // Expected: {'quot': 0, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 450,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b01010010; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 451,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00101100; // Expected: {'quot': 4, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 452,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b00000011; // Expected: {'quot': 75, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b00000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 453,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 75, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 454,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b00000110; // Expected: {'quot': 6, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 455,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 456,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b11001011; // Expected: {'quot': 0, 'rem': 119}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 457,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01000011; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 458,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10010110; // Expected: {'quot': 1, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 459,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b01011000; // Expected: {'quot': 0, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 460,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b00111101; // Expected: {'quot': 2, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 461,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 462,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 463,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01100111; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 464,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b00110100; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 465,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00110100; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 466,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 467,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b01001100; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 468,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 469,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b10011001; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 470,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 471,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 472,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01011100; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 473,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 474,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 475,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 476,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10000110; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 477,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01101001; // Expected: {'quot': 1, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 478,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 479,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01011010; // Expected: {'quot': 2, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 480,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b01011000; // Expected: {'quot': 2, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 481,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 482,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01110100; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 483,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b11001010; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 484,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10010111; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 485,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 177}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 486,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01010111; // Expected: {'quot': 2, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 487,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 206}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 488,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b01001000; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 489,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b11001001; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 490,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10000111; // Expected: {'quot': 1, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 491,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00101101; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 492,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 493,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10011110; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 494,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b01000000; // Expected: {'quot': 3, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 495,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 496,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00111101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 497,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 498,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 499,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00110001; // Expected: {'quot': 3, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 500,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00011100; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 501,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b11011011; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 502,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 503,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01001001; // Expected: {'quot': 2, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 504,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b01010011; // Expected: {'quot': 2, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 505,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00011110; // Expected: {'quot': 2, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 506,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 507,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 508,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b10011001; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 509,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b10010011; // Expected: {'quot': 0, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 510,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b00011011; // Expected: {'quot': 6, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 511,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 512,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10010001; // Expected: {'quot': 1, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 513,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 221}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 514,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 515,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00101000; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 516,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b01000000; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 517,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 518,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 519,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b10101110; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 520,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00011000; // Expected: {'quot': 3, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 521,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00010101; // Expected: {'quot': 5, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 522,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 523,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 524,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b01001000; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 525,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b01010101; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 526,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00001000; // Expected: {'quot': 18, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 527,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 18, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 528,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01000001; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 529,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 214}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 530,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 531,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00110011; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 532,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 533,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10100100; // Expected: {'quot': 1, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 534,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b00110010; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 535,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b00100111; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 536,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01111101; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 537,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b01101001; // Expected: {'quot': 2, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 538,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 539,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 540,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b01100010; // Expected: {'quot': 2, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 541,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b10010001; // Expected: {'quot': 0, 'rem': 133}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 542,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00010110; // Expected: {'quot': 3, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 543,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b01110111; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 544,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11100011; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 545,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b00101000; // Expected: {'quot': 1, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 546,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b01010111; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 547,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 548,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 549,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 550,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 551,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 552,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 553,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00010111; // Expected: {'quot': 7, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 554,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 555,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 556,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 557,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b00001010; // Expected: {'quot': 25, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 558,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 559,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 560,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b10100100; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b10100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 561,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 562,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b10001110; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 563,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 564,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00111111; // Expected: {'quot': 3, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 565,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 566,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b10110000; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 567,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b00001110; // Expected: {'quot': 16, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 568,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 16, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b01000001; // Expected: {'quot': 3, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 569,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01010110; // Expected: {'quot': 0, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 570,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 571,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b00001110; // Expected: {'quot': 11, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 572,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 127}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 573,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10101110; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 574,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b01000101; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 575,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 576,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01011001; // Expected: {'quot': 1, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 577,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 578,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b00000111; // Expected: {'quot': 24, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 579,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b01001001; // Expected: {'quot': 3, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 580,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 207}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 581,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00001101; // Expected: {'quot': 6, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 582,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b01001010; // Expected: {'quot': 3, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 583,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 584,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b01111010; // Expected: {'quot': 1, 'rem': 102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 585,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00111011; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 586,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 143}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 587,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11110100; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 588,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 589,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 590,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b00010100; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 591,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 592,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01111100; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 593,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 233}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 594,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b01110100; // Expected: {'quot': 1, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 595,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b01011011; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 596,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b01010011; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 597,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b00101000; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 598,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 599,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00100001; // Expected: {'quot': 4, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 600,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01101011; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 601,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b01111001; // Expected: {'quot': 1, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 602,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b11010001; // Expected: {'quot': 1, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 603,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b01110111; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 604,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01101010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 605,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b11110011; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b11110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 606,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01000110; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 607,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00101010; // Expected: {'quot': 5, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 608,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b00001110; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 609,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00000101; // Expected: {'quot': 43, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 610,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 43, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 611,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 612,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b00110010; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 613,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b00110010; // Expected: {'quot': 3, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 614,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b00110010; // Expected: {'quot': 2, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 615,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 616,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b01010010; // Expected: {'quot': 2, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 617,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b10111111; // Expected: {'quot': 1, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 618,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 619,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 620,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00101110; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 621,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b00110101; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b00110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 622,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b11001101; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 623,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 624,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 625,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01100001; // Expected: {'quot': 1, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 626,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 627,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01101110; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 628,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01111010; // Expected: {'quot': 1, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 629,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00010000; // Expected: {'quot': 15, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 630,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b10100000; // Expected: {'quot': 1, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 631,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b00000100; // Expected: {'quot': 17, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b00000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 632,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b01101110; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 633,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10011110; // Expected: {'quot': 0, 'rem': 149}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 634,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01010011; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 635,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00011111; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 636,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 637,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 638,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10001000; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 639,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 640,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b00000010; // Expected: {'quot': 90, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 641,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 90, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b01011001; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 642,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b01100101; // Expected: {'quot': 2, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 643,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 644,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b01011110; // Expected: {'quot': 0, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b01011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 645,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 646,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 647,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b11000101; // Expected: {'quot': 0, 'rem': 159}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 648,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01011111; // Expected: {'quot': 1, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 649,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01001000; // Expected: {'quot': 2, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 650,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b10000010; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 651,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 652,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 653,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00100111; // Expected: {'quot': 5, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 654,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 655,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b00101010; // Expected: {'quot': 3, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 656,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b11011000; // Expected: {'quot': 0, 'rem': 210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 657,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00000011; // Expected: {'quot': 64, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 658,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 64, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00101110; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 659,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10011100; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 660,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b01101000; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 661,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01101000; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 662,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b10000000; // Expected: {'quot': 1, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 663,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10100010; // Expected: {'quot': 0, 'rem': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 664,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 665,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00011000; // Expected: {'quot': 8, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 666,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10101001; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 667,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 668,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b00101100; // Expected: {'quot': 3, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 669,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 670,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01001001; // Expected: {'quot': 3, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 671,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 672,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01001110; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 673,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b00011111; // Expected: {'quot': 2, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 674,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b01100110; // Expected: {'quot': 2, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 675,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10111100; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 676,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01011101; // Expected: {'quot': 2, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 677,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b01100111; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 678,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 679,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b01110001; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 680,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01011011; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 681,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10100110; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 682,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 683,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01000001; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 684,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 685,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00111111; // Expected: {'quot': 3, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 686,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b00001000; // Expected: {'quot': 27, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 687,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 27, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b01111111; // Expected: {'quot': 1, 'rem': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 688,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01000110; // Expected: {'quot': 3, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 689,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b10110100; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 690,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 213}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 691,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 692,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 693,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b10000010; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 694,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b01001000; // Expected: {'quot': 2, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 695,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 696,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b01101000; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 697,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b01011111; // Expected: {'quot': 0, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 698,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 699,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 700,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b00110001; // Expected: {'quot': 3, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 701,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01100100; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 702,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b01011000; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 703,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 704,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b00101110; // Expected: {'quot': 4, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 705,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b01010010; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 706,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 707,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10000011; // Expected: {'quot': 1, 'rem': 102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 708,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b10101001; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 709,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 710,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00110001; // Expected: {'quot': 4, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 711,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01101110; // Expected: {'quot': 1, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 712,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b00100101; // Expected: {'quot': 6, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 713,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00111000; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 714,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 715,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 716,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 717,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01011010; // Expected: {'quot': 2, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 718,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00001011; // Expected: {'quot': 17, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 719,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 720,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b00101011; // Expected: {'quot': 5, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 721,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 722,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00101000; // Expected: {'quot': 4, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 723,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00110110; // Expected: {'quot': 3, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 724,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10010010; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 725,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10101110; // Expected: {'quot': 1, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 726,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b01001111; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 727,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 728,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01000010; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 729,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 730,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 731,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b00000101; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 732,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11010011; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 733,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 734,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01010110; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 735,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 157}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 736,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 191}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 737,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b00111010; // Expected: {'quot': 1, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 738,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 739,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00100010; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 740,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 741,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b00010110; // Expected: {'quot': 7, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 742,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b10001000; // Expected: {'quot': 1, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 743,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b10000010; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 744,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 745,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b11001101; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 746,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 747,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b10001101; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 748,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b00011010; // Expected: {'quot': 3, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 749,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10001000; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 750,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 751,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01001100; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 752,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 753,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b00010000; // Expected: {'quot': 15, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 754,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 755,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00101100; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 756,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 188}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 757,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b10011111; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 758,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 759,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01000111; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 760,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b01101011; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 761,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b11000100; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 762,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b11011000; // Expected: {'quot': 0, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 763,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b10010101; // Expected: {'quot': 1, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b10010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 764,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b01100010; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 765,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00101011; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 766,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 767,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b10110011; // Expected: {'quot': 0, 'rem': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 768,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 769,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00000001; // Expected: {'quot': 63, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 770,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00001010; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 771,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b11001010; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 772,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 773,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10100011; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 774,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 775,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b00101000; // Expected: {'quot': 4, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 776,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01000111; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 777,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00100010; // Expected: {'quot': 5, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 778,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 779,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 780,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 781,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b00000111; // Expected: {'quot': 19, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 782,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 19, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 783,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b01100011; // Expected: {'quot': 2, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 784,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00010011; // Expected: {'quot': 9, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 785,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b10000101; // Expected: {'quot': 0, 'rem': 130}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 786,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b00101001; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 787,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b01101001; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 788,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 789,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 790,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11011001; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 791,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 792,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b00100001; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 793,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11110011; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 794,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b10001111; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 795,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 796,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10101111; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 797,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b01011001; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 798,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b10000111; // Expected: {'quot': 1, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 799,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b00110100; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 800,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 801,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10000101; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 802,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b00100101; // Expected: {'quot': 2, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 803,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 804,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 805,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b10011110; // Expected: {'quot': 0, 'rem': 157}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 806,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10110001; // Expected: {'quot': 1, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 807,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00011100; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 808,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b01001111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 809,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 810,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 811,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 169}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 812,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 813,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 814,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11010011; // Expected: {'quot': 0, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 815,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 816,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b00111100; // Expected: {'quot': 2, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 817,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b01011110; // Expected: {'quot': 2, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b01011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 818,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01011011; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 819,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 820,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11101011; // Expected: {'quot': 0, 'rem': 142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 821,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 822,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b00101010; // Expected: {'quot': 5, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 823,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01001000; // Expected: {'quot': 2, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 824,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b00001101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 825,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 826,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10111011; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 827,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b10100010; // Expected: {'quot': 0, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 828,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 829,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00000010; // Expected: {'quot': 61, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 830,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 61, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 831,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 832,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b00011001; // Expected: {'quot': 9, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b00011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 833,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00111010; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 834,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b11010010; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 835,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00011000; // Expected: {'quot': 7, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 836,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01100010; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 837,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 838,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10101001; // Expected: {'quot': 1, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 839,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 840,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 157}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 841,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11000101; // Expected: {'quot': 0, 'rem': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 842,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 843,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 844,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b00111101; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 845,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b11000000; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 846,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b00111011; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 847,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b00001111; // Expected: {'quot': 4, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 848,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 849,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00011111; // Expected: {'quot': 3, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 850,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10111011; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 851,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01110001; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 852,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00010011; // Expected: {'quot': 9, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 853,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b00001101; // Expected: {'quot': 3, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 854,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01001101; // Expected: {'quot': 1, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 855,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 134}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 856,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b00001100; // Expected: {'quot': 16, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 857,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 16, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b01011010; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 858,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b10111010; // Expected: {'quot': 1, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 859,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 860,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00010001; // Expected: {'quot': 5, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 861,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b01111011; // Expected: {'quot': 1, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 862,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 863,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b01011111; // Expected: {'quot': 2, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 864,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b01000000; // Expected: {'quot': 3, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 865,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b00100111; // Expected: {'quot': 6, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 866,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10101000; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 867,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00000010; // Expected: {'quot': 24, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 868,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 24, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01101110; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 869,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 870,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 871,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b00010111; // Expected: {'quot': 9, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 872,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01011111; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 873,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 874,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b10001001; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 875,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 876,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 877,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 878,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b10111011; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 879,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01000010; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 880,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 881,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 882,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b00100010; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 883,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b00011101; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b00011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 884,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 885,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10110010; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 886,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 887,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 888,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b00110100; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 889,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 890,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10000100; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 891,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b01001101; // Expected: {'quot': 3, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 892,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 893,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b00001011; // Expected: {'quot': 13, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 894,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00011110; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 895,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00010001; // Expected: {'quot': 10, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 896,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00011111; // Expected: {'quot': 3, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 897,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01110100; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 898,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 899,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 900,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 115}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 901,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 902,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 903,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 904,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b10001000; // Expected: {'quot': 1, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 905,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10010111; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 906,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b00101111; // Expected: {'quot': 3, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 907,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b10001011; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 908,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00101111; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 909,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b00011110; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 910,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00100100; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 911,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 912,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 913,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b10001001; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 914,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 915,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10011110; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 916,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b01101100; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b01101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 917,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01001100; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 918,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b11010111; // Expected: {'quot': 1, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 919,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b00011010; // Expected: {'quot': 4, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 920,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 921,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 922,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b11101011; // Expected: {'quot': 0, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 923,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b01101100; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b01101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 924,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 925,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b00110011; // Expected: {'quot': 3, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 926,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01000011; // Expected: {'quot': 2, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 927,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b01011010; // Expected: {'quot': 1, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 928,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00001101; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 929,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 930,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 931,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 932,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 933,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00111111; // Expected: {'quot': 3, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 934,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b01011001; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 935,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 936,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 937,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00001010; // Expected: {'quot': 12, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 938,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b10001011; // Expected: {'quot': 1, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 939,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 940,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 941,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 942,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b01111001; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 943,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b00010001; // Expected: {'quot': 10, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 944,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b00010111; // Expected: {'quot': 6, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 945,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b00101011; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 946,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01111100; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 947,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b00111001; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 948,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00001000; // Expected: {'quot': 25, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 949,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b01000000; // Expected: {'quot': 2, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 950,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b01000001; // Expected: {'quot': 1, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 951,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01101010; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 952,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 953,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b01000011; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 954,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b00000001; // Expected: {'quot': 195, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 955,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 195, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b10001010; // Expected: {'quot': 0, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 956,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b00001111; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 957,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b10011110; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 958,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 959,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b10100000; // Expected: {'quot': 0, 'rem': 115}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 960,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b10010001; // Expected: {'quot': 1, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 961,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 962,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b01100101; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 963,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b00101001; // Expected: {'quot': 5, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 964,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 965,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b01011100; // Expected: {'quot': 0, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 966,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b10000001; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 967,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b00110101; // Expected: {'quot': 2, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b00110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 968,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b00111110; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 969,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01101010; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 970,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b11100111; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 971,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b01010000; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 972,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00110011; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 973,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b11100010; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 974,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b01100101; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 975,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b00010100; // Expected: {'quot': 6, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 976,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b01011110; // Expected: {'quot': 0, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b01011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 977,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 978,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 979,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b00010001; // Expected: {'quot': 12, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 980,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 981,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 982,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b01000110; // Expected: {'quot': 2, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 983,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b01110100; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 984,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b11010101; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 985,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01100001; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 986,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 987,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b00111101; // Expected: {'quot': 3, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 988,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b10000101; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 989,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 990,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00111100; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 991,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 992,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 993,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b00000110; // Expected: {'quot': 35, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 994,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 35, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b11001101; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 995,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b11011011; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 996,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 997,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b00110110; // Expected: {'quot': 4, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 998,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b00000010; // Expected: {'quot': 109, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 999,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 109, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b10001000; // Expected: {'quot': 1, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1000,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1001,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b10001110; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1002,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 109}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1003,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00111011; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1004,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1005,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b00110100; // Expected: {'quot': 2, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1006,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b00000011; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b00000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1007,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b00111001; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1008,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01000111; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1009,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11000110; // Expected: {'quot': 1, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1010,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1011,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 248}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1012,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1013,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1014,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1015,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 149}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1016,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01100010; // Expected: {'quot': 1, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1017,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1018,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b10100110; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b10100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1019,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b01110000; // Expected: {'quot': 1, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1020,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b00111000; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1021,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00010110; // Expected: {'quot': 5, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1022,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1023,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1024,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01000010; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1025,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10011101; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1026,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10100011; // Expected: {'quot': 1, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1027,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11001010; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1028,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00101010; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1029,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00011010; // Expected: {'quot': 4, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1030,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b10100011; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1031,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b01010110; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1032,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10110010; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1033,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b01001001; // Expected: {'quot': 2, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1034,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1035,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1036,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1037,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b00101110; // Expected: {'quot': 3, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1038,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00111100; // Expected: {'quot': 3, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1039,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 161}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1040,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01100001; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1041,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1042,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1043,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01011111; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1044,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00011011; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1045,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b10001100; // Expected: {'quot': 1, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1046,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01110111; // Expected: {'quot': 2, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1047,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1048,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b00011101; // Expected: {'quot': 8, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b00011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1049,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b00101000; // Expected: {'quot': 4, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1050,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01101000; // Expected: {'quot': 1, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1051,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1052,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b00000110; // Expected: {'quot': 36, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1053,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 36, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b10001010; // Expected: {'quot': 0, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1054,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b01000001; // Expected: {'quot': 2, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1055,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1056,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10000100; // Expected: {'quot': 1, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1057,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b00001101; // Expected: {'quot': 12, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1058,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b00110100; // Expected: {'quot': 4, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1059,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1060,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1061,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b01111001; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1062,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b11001010; // Expected: {'quot': 0, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1063,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b00110000; // Expected: {'quot': 4, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1064,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b00101101; // Expected: {'quot': 5, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1065,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01011011; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1066,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b01010100; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1067,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1068,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1069,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 191}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1070,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1071,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b00010101; // Expected: {'quot': 8, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1072,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1073,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 222}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1074,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11101011; // Expected: {'quot': 0, 'rem': 217}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1075,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10000010; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1076,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b00010011; // Expected: {'quot': 10, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1077,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1078,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b10101111; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1079,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01110100; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1080,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01110001; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1081,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01000001; // Expected: {'quot': 2, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1082,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b10011010; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1083,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01110000; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1084,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00110000; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1085,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1086,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11000110; // Expected: {'quot': 1, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1087,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b01111011; // Expected: {'quot': 1, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1088,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b01000101; // Expected: {'quot': 2, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1089,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10001010; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1090,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01011001; // Expected: {'quot': 2, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1091,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b01111111; // Expected: {'quot': 1, 'rem': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1092,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1093,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01101110; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1094,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1095,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1096,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1097,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b01000000; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1098,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00110000; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1099,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00111010; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1100,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10100000; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1101,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 202}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1102,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1103,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b10001100; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1104,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b01000000; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1105,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b00100011; // Expected: {'quot': 4, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1106,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1107,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00101011; // Expected: {'quot': 4, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1108,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 202}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1109,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00111110; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1110,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11001000; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1111,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11001010; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1112,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b10000101; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1113,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b00001010; // Expected: {'quot': 14, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1114,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b00010010; // Expected: {'quot': 12, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b00010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1115,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1116,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b01011000; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1117,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1118,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1119,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b10100011; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1120,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b01100101; // Expected: {'quot': 2, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1121,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b00000010; // Expected: {'quot': 93, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1122,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 93, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b00101000; // Expected: {'quot': 5, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1123,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b10000000; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1124,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b00011101; // Expected: {'quot': 5, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b00011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1125,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1126,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b00111111; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1127,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b00001110; // Expected: {'quot': 14, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1128,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1129,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10010100; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1130,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1131,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00000001; // Expected: {'quot': 249, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1132,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 249, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b00010101; // Expected: {'quot': 8, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1133,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00111111; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1134,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b00101010; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1135,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b00101101; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1136,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b00001010; // Expected: {'quot': 8, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1137,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01000100; // Expected: {'quot': 2, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1138,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1139,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1140,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00011110; // Expected: {'quot': 3, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1141,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b00111100; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1142,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1143,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b01100001; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1144,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b00101111; // Expected: {'quot': 1, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1145,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10000010; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1146,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b00000010; // Expected: {'quot': 38, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1147,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 38, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b00010100; // Expected: {'quot': 2, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1148,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00001001; // Expected: {'quot': 26, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1149,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 26, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00111100; // Expected: {'quot': 2, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1150,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00011000; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1151,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b01000110; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1152,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b00001001; // Expected: {'quot': 25, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b00001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1153,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 25, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1154,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01111000; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1155,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1156,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1157,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00101100; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1158,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01000111; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1159,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01010001; // Expected: {'quot': 1, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1160,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1161,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b01001001; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1162,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1163,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 179}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1164,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1165,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00001001; // Expected: {'quot': 16, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1166,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 16, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1167,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00010000; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1168,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01100110; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1169,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b01011100; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1170,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1171,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 181}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1172,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 163}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1173,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01011000; // Expected: {'quot': 1, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1174,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10110000; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1175,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b00011010; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1176,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b00000110; // Expected: {'quot': 26, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1177,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 26, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b00101111; // Expected: {'quot': 4, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1178,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1179,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b10100101; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1180,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b01110011; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1181,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b01000101; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1182,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 180}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1183,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b00001100; // Expected: {'quot': 10, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1184,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1185,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b10001101; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1186,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10111000; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1187,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11010100; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1188,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1189,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00001010; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1190,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00010001; // Expected: {'quot': 11, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1191,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11011111; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1192,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1193,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1194,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1195,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b11110011; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b11110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1196,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1197,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01101000; // Expected: {'quot': 0, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1198,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1199,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b01011101; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1200,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01100101; // Expected: {'quot': 1, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1201,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b01100100; // Expected: {'quot': 0, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1202,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b10000110; // Expected: {'quot': 0, 'rem': 119}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1203,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b11000100; // Expected: {'quot': 1, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1204,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1205,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b10101001; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1206,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00110101; // Expected: {'quot': 3, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1207,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10110101; // Expected: {'quot': 1, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1208,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b10111001; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1209,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b10110100; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1210,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b01100000; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1211,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1212,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1213,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1214,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1215,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00011010; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1216,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b01110100; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1217,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b00010111; // Expected: {'quot': 5, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1218,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10011111; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1219,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01100111; // Expected: {'quot': 2, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1220,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b00110010; // Expected: {'quot': 2, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1221,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10001101; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1222,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b00111000; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1223,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11000011; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1224,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b10101100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1225,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10101110; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1226,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00001011; // Expected: {'quot': 14, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1227,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1228,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b01000111; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1229,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b01010100; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1230,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b01001100; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1231,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01100110; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1232,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1233,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b10100011; // Expected: {'quot': 0, 'rem': 114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1234,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00000110; // Expected: {'quot': 41, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1235,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 41, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1236,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b00001010; // Expected: {'quot': 12, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1237,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1238,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1239,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00111100; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1240,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01101100; // Expected: {'quot': 1, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1241,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 151}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1242,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b00000111; // Expected: {'quot': 27, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1243,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 27, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b01110001; // Expected: {'quot': 0, 'rem': 111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1244,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01101010; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1245,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1246,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1247,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1248,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b10110011; // Expected: {'quot': 0, 'rem': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1249,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01100111; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1250,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b10011000; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1251,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b10000000; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1252,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b01111111; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1253,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10110100; // Expected: {'quot': 0, 'rem': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1254,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01001101; // Expected: {'quot': 1, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1255,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111100; Y = 8'b01111110; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111100; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1256,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1257,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b00101101; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1258,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b10110100; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1259,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1260,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00010100; // Expected: {'quot': 9, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1261,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b01011011; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1262,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b11001001; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1263,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b01010110; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1264,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b01110000; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1265,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01000100; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1266,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b00100000; // Expected: {'quot': 4, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b00100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1267,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10110000; // Expected: {'quot': 1, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1268,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00001010; // Expected: {'quot': 8, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1269,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00010110; // Expected: {'quot': 9, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1270,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b10001111; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1271,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b00010000; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1272,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b10101100; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1273,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 210}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1274,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1275,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1276,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00101100; // Expected: {'quot': 3, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1277,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1278,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1279,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b01011100; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1280,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1281,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1282,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01101100; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1283,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b00110000; // Expected: {'quot': 3, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1284,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000010; Y = 8'b00101010; // Expected: {'quot': 3, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000010; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1285,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b00110110; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1286,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1287,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01101010; // Expected: {'quot': 2, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1288,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b00000101; // Expected: {'quot': 42, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1289,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 42, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01010101; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1290,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10101000; // Expected: {'quot': 1, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1291,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b01101111; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1292,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b00000111; // Expected: {'quot': 17, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1293,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00011001; // Expected: {'quot': 4, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1294,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b01001110; // Expected: {'quot': 2, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1295,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1296,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b01100100; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1297,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b00010111; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1298,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b00100110; // Expected: {'quot': 5, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b00100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1299,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b00110110; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1300,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1301,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b10010100; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1302,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10110011; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1303,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10010011; // Expected: {'quot': 1, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1304,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b00111010; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1305,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1306,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1307,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01001010; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1308,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b10111000; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1309,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b00111110; // Expected: {'quot': 3, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1310,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b10011010; // Expected: {'quot': 0, 'rem': 139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1311,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01101110; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1312,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1313,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00110000; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1314,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b10010001; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1315,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b00100010; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1316,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01101101; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1317,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 241}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1318,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1319,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10000001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1320,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01010111; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1321,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10100000; // Expected: {'quot': 1, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1322,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b11001001; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1323,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1324,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01110001; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1325,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b01111111; // Expected: {'quot': 1, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1326,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10100111; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1327,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b10010001; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1328,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b00001110; // Expected: {'quot': 3, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1329,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00101001; // Expected: {'quot': 5, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1330,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10111111; // Expected: {'quot': 1, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1331,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b00110100; // Expected: {'quot': 3, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1332,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b11011110; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1333,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b00101111; // Expected: {'quot': 3, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1334,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11000000; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1335,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110010; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110010; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1336,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01101101; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1337,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b11000110; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1338,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b10001011; // Expected: {'quot': 1, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1339,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11011000; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1340,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1341,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b01001111; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1342,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b00010111; // Expected: {'quot': 5, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1343,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b01010100; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1344,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01100100; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1345,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00011110; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1346,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b10101010; // Expected: {'quot': 1, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1347,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1348,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1349,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b10110111; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1350,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1351,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b10100010; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1352,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b00101011; // Expected: {'quot': 3, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1353,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1354,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1355,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1356,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b01010011; // Expected: {'quot': 0, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1357,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b00000001; // Expected: {'quot': 66, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1358,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 66, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b00101010; // Expected: {'quot': 3, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1359,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00001110; // Expected: {'quot': 17, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1360,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b00001010; // Expected: {'quot': 15, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1361,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b10110000; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1362,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1363,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1364,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b00101000; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1365,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b01111001; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1366,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1367,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b01100111; // Expected: {'quot': 2, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1368,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1369,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1370,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b00110001; // Expected: {'quot': 3, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1371,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b00010011; // Expected: {'quot': 8, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1372,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b00101101; // Expected: {'quot': 3, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1373,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1374,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b00100101; // Expected: {'quot': 5, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1375,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00010000; // Expected: {'quot': 8, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1376,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 115}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1377,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b10010101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b10010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1378,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00011010; // Expected: {'quot': 9, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1379,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b00101101; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1380,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00111010; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1381,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1382,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b00011010; // Expected: {'quot': 6, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1383,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b01011010; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1384,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1385,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00111011; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1386,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1387,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b01101101; // Expected: {'quot': 0, 'rem': 102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b01101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1388,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b00001010; // Expected: {'quot': 16, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1389,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 16, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b00010001; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1390,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00111101; // Expected: {'quot': 3, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1391,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01100010; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1392,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01101001; // Expected: {'quot': 1, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1393,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1394,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1395,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1396,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b00001110; // Expected: {'quot': 14, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1397,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01110000; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1398,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b10000001; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1399,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1400,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b00000110; // Expected: {'quot': 36, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1401,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 36, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b10000111; // Expected: {'quot': 1, 'rem': 114}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1402,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1403,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b11010011; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1404,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b10011110; // Expected: {'quot': 0, 'rem': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1405,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b01000100; // Expected: {'quot': 3, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1406,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b00011111; // Expected: {'quot': 5, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1407,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1408,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b11101100; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1409,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01001110; // Expected: {'quot': 1, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1410,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b01010000; // Expected: {'quot': 2, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1411,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b10101100; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1412,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1413,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b01011110; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b01011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1414,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b01011010; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1415,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b11111010; // Expected: {'quot': 0, 'rem': 163}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1416,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1417,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b01001110; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1418,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1419,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1420,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b11000111; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1421,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00010001; // Expected: {'quot': 6, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1422,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00001010; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1423,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b00110010; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1424,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b01010101; // Expected: {'quot': 3, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1425,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00011000; // Expected: {'quot': 7, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1426,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b10000010; // Expected: {'quot': 0, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1427,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01011010; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1428,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1429,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b00100010; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1430,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b01000001; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1431,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00001011; // Expected: {'quot': 11, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1432,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00001110; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1433,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1434,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01000011; // Expected: {'quot': 2, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1435,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1436,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b01011100; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1437,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 143}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1438,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01001110; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1439,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b11001011; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1440,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01111010; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1441,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b00011111; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1442,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b10001101; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1443,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00111010; // Expected: {'quot': 4, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1444,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1445,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b00111101; // Expected: {'quot': 3, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1446,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 123}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1447,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1448,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00110101; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1449,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b01010010; // Expected: {'quot': 2, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1450,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1451,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10001010; // Expected: {'quot': 1, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1452,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00001100; // Expected: {'quot': 8, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1453,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b01001100; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1454,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01110010; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1455,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1456,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1457,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b01100001; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1458,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01000011; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1459,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1460,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b01000000; // Expected: {'quot': 3, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1461,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1462,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01111111; // Expected: {'quot': 0, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1463,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b01100001; // Expected: {'quot': 1, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1464,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1465,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b01011101; // Expected: {'quot': 2, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1466,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1467,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b01111111; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1468,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10100001; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1469,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b10101001; // Expected: {'quot': 1, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1470,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1471,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10101101; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1472,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1473,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b00100111; // Expected: {'quot': 2, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1474,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10010000; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1475,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b01010000; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1476,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b01100001; // Expected: {'quot': 1, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1477,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10010010; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1478,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00000101; // Expected: {'quot': 29, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1479,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 29, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b00110010; // Expected: {'quot': 4, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1480,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1481,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1482,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01100000; // Expected: {'quot': 1, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1483,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1484,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00100110; // Expected: {'quot': 5, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1485,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01111010; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1486,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00010100; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1487,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1488,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1489,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1490,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b00110001; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1491,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b10000010; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1492,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1493,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b10101111; // Expected: {'quot': 1, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1494,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1495,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1496,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1497,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01111010; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1498,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b00001010; // Expected: {'quot': 9, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1499,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1500,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1501,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1502,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10001000; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1503,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1504,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1505,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 202}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1506,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1507,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10101001; // Expected: {'quot': 1, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1508,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b01101001; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1509,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b10001100; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1510,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1511,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1512,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11001011; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1513,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 163}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1514,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1515,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 163}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1516,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b01101001; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1517,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b01110011; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1518,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b01010010; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1519,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1520,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 149}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1521,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b01000111; // Expected: {'quot': 3, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1522,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1523,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1524,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01110100; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1525,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00010001; // Expected: {'quot': 4, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1526,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01001010; // Expected: {'quot': 1, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1527,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b01100111; // Expected: {'quot': 1, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1528,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1529,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b00101011; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1530,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1531,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b11100011; // Expected: {'quot': 0, 'rem': 178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1532,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1533,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1534,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b01000100; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1535,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 191}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1536,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1537,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b00011110; // Expected: {'quot': 4, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1538,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1539,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010000; Y = 8'b00100110; // Expected: {'quot': 5, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010000; Y = 8'b00100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1540,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b00010110; // Expected: {'quot': 3, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1541,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01011001; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1542,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1543,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1544,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00011010; // Expected: {'quot': 6, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1545,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1546,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10001010; // Expected: {'quot': 1, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1547,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1548,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b01100111; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1549,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b10010110; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1550,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1551,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1552,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10100010; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1553,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b11011100; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1554,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01111100; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1555,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b01110001; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1556,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1557,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1558,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b00110100; // Expected: {'quot': 3, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1559,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b10011111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1560,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00111100; // Expected: {'quot': 2, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1561,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1562,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11001001; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1563,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1564,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00010101; // Expected: {'quot': 11, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1565,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1566,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10011101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1567,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b00110110; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1568,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b01000100; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1569,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01110011; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1570,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1571,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b00100111; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1572,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1573,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1574,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b00011001; // Expected: {'quot': 6, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b00011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1575,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10010001; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1576,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b01100100; // Expected: {'quot': 1, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1577,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b10100000; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1578,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1579,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00101001; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1580,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11001011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1581,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b00010010; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b00010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1582,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1583,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b00100010; // Expected: {'quot': 5, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1584,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00010100; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1585,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1586,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b00100101; // Expected: {'quot': 3, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1587,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01111000; // Expected: {'quot': 1, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1588,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11001111; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1589,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1590,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1591,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1592,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1593,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100001; Y = 8'b00100011; // Expected: {'quot': 4, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100001; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1594,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101101; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 173}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101101; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1595,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1596,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00000110; // Expected: {'quot': 26, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1597,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 26, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1598,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1599,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1600,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 175}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1601,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00001101; // Expected: {'quot': 18, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1602,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 18, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00011100; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1603,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b10110001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1604,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b11010011; // Expected: {'quot': 0, 'rem': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1605,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b01001100; // Expected: {'quot': 2, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1606,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b10010111; // Expected: {'quot': 0, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1607,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 202}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1608,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1609,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b10110111; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1610,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1611,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1612,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b11001000; // Expected: {'quot': 1, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1613,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1614,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 226}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1615,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11001011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1616,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00010001; // Expected: {'quot': 7, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1617,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1618,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b00100010; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1619,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1620,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00011100; // Expected: {'quot': 7, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1621,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1622,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1623,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b00001011; // Expected: {'quot': 9, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1624,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1625,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b01101101; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b01101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1626,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b01001000; // Expected: {'quot': 2, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1627,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1628,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01100111; // Expected: {'quot': 1, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1629,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01111000; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1630,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01011001; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1631,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1632,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b01001000; // Expected: {'quot': 3, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1633,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11001011; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1634,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b00001001; // Expected: {'quot': 13, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b00001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1635,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b11000101; // Expected: {'quot': 0, 'rem': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1636,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b00101011; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1637,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1638,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b01001111; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1639,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1640,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00100000; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1641,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 169}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1642,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b10111101; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1643,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10111101; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1644,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 119}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1645,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10111010; // Expected: {'quot': 1, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1646,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 181}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1647,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00001000; // Expected: {'quot': 31, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1648,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 31, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b10011111; // Expected: {'quot': 0, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1649,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b10110111; // Expected: {'quot': 0, 'rem': 125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1650,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1651,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1652,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1653,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01011100; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1654,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b01011110; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b01011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1655,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1656,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 116}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1657,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b00010100; // Expected: {'quot': 6, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1658,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1659,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b10111111; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1660,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01000100; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1661,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1662,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b00011110; // Expected: {'quot': 4, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1663,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01111100; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1664,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1665,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b00010100; // Expected: {'quot': 3, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1666,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1667,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1668,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01100100; // Expected: {'quot': 0, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1669,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 112}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1670,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b00100111; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1671,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 169}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1672,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01111000; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1673,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b10111111; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1674,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b10011010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1675,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1676,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b00101001; // Expected: {'quot': 4, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1677,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 149}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1678,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b01111110; // Expected: {'quot': 1, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1679,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b10010001; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1680,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00001010; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1681,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1682,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b00011011; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1683,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1684,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1685,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 137}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1686,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10001101; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1687,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b00110010; // Expected: {'quot': 4, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1688,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00101000; // Expected: {'quot': 3, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1689,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01011000; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1690,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b01001000; // Expected: {'quot': 3, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1691,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00110110; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1692,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1693,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b00110010; // Expected: {'quot': 3, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1694,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1695,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1696,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b10100010; // Expected: {'quot': 0, 'rem': 148}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1697,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110011; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 115}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110011; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1698,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10100010; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1699,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10101111; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1700,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10001100; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1701,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b00110111; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b00110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1702,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01001000; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1703,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1704,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10111000; // Expected: {'quot': 0, 'rem': 169}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1705,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b00011000; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1706,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b10000111; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1707,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1708,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b10000001; // Expected: {'quot': 1, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1709,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10101011; // Expected: {'quot': 1, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1710,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1711,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b00001011; // Expected: {'quot': 5, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1712,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 167}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1713,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b00111011; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1714,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b01000110; // Expected: {'quot': 3, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1715,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00111100; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1716,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1717,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1718,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 233}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1719,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b00011111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1720,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b10100010; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1721,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b01010111; // Expected: {'quot': 2, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1722,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b11010001; // Expected: {'quot': 0, 'rem': 181}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b11010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1723,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01011101; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1724,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01000100; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1725,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01111100; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1726,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b00001100; // Expected: {'quot': 17, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1727,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1728,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b00011001; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b00011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1729,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00111010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1730,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1731,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1732,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10011101; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1733,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10000010; // Expected: {'quot': 1, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1734,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b00101110; // Expected: {'quot': 3, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1735,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011100; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 92}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011100; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1736,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00110111; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1737,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11011111; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1738,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b00110101; // Expected: {'quot': 3, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b00110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1739,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00101101; // Expected: {'quot': 2, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1740,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b00000111; // Expected: {'quot': 29, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1741,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 29, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1742,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b01001000; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1743,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b01001111; // Expected: {'quot': 1, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1744,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b00011110; // Expected: {'quot': 6, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1745,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1746,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b01010111; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1747,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00110011; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1748,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1749,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b00011000; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1750,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00100110; // Expected: {'quot': 5, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1751,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10100100; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1752,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1753,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b01001111; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1754,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b01011000; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1755,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00010010; // Expected: {'quot': 7, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1756,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b01010110; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1757,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b01101011; // Expected: {'quot': 1, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1758,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1759,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11010110; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1760,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b00100100; // Expected: {'quot': 4, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1761,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01011010; // Expected: {'quot': 1, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1762,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1763,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10001000; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1764,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 182}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1765,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01010001; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1766,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b11100011; // Expected: {'quot': 0, 'rem': 145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1767,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b01111101; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b01111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1768,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10000111; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1769,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b00101101; // Expected: {'quot': 4, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1770,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b01101100; // Expected: {'quot': 0, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b01101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1771,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b01001110; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1772,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1773,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b00100111; // Expected: {'quot': 1, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1774,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10100100; // Expected: {'quot': 0, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1775,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b00100100; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1776,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b10001111; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1777,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1778,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b10011011; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1779,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10000101; // Expected: {'quot': 1, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1780,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1781,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1782,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10011111; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1783,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b00111111; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1784,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b00111111; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1785,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b00010010; // Expected: {'quot': 7, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b00010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1786,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b10101011; // Expected: {'quot': 0, 'rem': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b10101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1787,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00010011; // Expected: {'quot': 12, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1788,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1789,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1790,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00111011; // Expected: {'quot': 1, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1791,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1792,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b01101011; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1793,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01001010; // Expected: {'quot': 1, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1794,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1795,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1796,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1797,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1798,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b01000111; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1799,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b01000010; // Expected: {'quot': 2, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1800,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11101100; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1801,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1802,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1803,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1804,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b00110010; // Expected: {'quot': 4, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1805,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b00110111; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b00110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1806,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00111101; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1807,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10101101; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1808,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b00011011; // Expected: {'quot': 2, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1809,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b00010110; // Expected: {'quot': 8, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1810,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01101101; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1811,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b00010011; // Expected: {'quot': 8, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1812,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00100010; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1813,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b10101000; // Expected: {'quot': 1, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1814,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 191}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1815,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b00010111; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1816,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b00011110; // Expected: {'quot': 5, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1817,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10100011; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1818,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00100010; // Expected: {'quot': 7, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1819,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00110000; // Expected: {'quot': 2, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1820,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b10011111; // Expected: {'quot': 0, 'rem': 145}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1821,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00001010; // Expected: {'quot': 8, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1822,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b00111100; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1823,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b00111110; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1824,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1825,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001001; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 201}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001001; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1826,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b01100101; // Expected: {'quot': 2, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1827,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1828,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b01011011; // Expected: {'quot': 2, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1829,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00100001; // Expected: {'quot': 2, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1830,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 207}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1831,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01001001; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1832,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b01110100; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1833,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01100110; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1834,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b01101110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1835,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b10111111; // Expected: {'quot': 0, 'rem': 185}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1836,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b11101011; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1837,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b10010111; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1838,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10010100; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1839,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b01000011; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1840,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1841,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b00010100; // Expected: {'quot': 9, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1842,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b01100001; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1843,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1844,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11000100; // Expected: {'quot': 1, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1845,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1846,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b00011110; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1847,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b11100011; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1848,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1849,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b10011111; // Expected: {'quot': 1, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1850,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1851,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b00011010; // Expected: {'quot': 8, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1852,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01110000; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1853,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b10100000; // Expected: {'quot': 0, 'rem': 154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1854,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1855,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 176}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1856,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01101010; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1857,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01001110; // Expected: {'quot': 2, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1858,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b00001111; // Expected: {'quot': 4, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1859,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b01010001; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b01010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1860,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10110011; // Expected: {'quot': 0, 'rem': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1861,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001101; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001101; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1862,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1863,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b01111001; // Expected: {'quot': 0, 'rem': 96}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1864,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01001101; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1865,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10111011; // Expected: {'quot': 0, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1866,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b00001011; // Expected: {'quot': 6, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1867,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1868,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b10011111; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1869,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00001101; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1870,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00100111; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1871,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1872,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b00110010; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1873,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00100000; // Expected: {'quot': 5, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1874,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b01111110; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1875,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b01010110; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1876,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b01101111; // Expected: {'quot': 1, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b01101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1877,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b00011100; // Expected: {'quot': 4, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1878,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01110010; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1879,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00001101; // Expected: {'quot': 16, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1880,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 16, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b01000111; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1881,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1882,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b11001001; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1883,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1884,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00010001; // Expected: {'quot': 14, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1885,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1886,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1887,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b10100101; // Expected: {'quot': 1, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1888,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b01110000; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1889,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1890,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b01000011; // Expected: {'quot': 1, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1891,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b01001110; // Expected: {'quot': 2, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1892,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01010101; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1893,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b00110011; // Expected: {'quot': 1, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1894,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b01101001; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1895,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b00110111; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b00110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1896,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1897,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b00011011; // Expected: {'quot': 5, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1898,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1899,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b11000111; // Expected: {'quot': 0, 'rem': 184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b11000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1900,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b11100011; // Expected: {'quot': 0, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1901,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1902,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1903,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b00110100; // Expected: {'quot': 4, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1904,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10011000; // Expected: {'quot': 1, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1905,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1906,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1907,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1908,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00100101; // Expected: {'quot': 3, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1909,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b11000110; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1910,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1911,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00101011; // Expected: {'quot': 1, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1912,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000011; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000011; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1913,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1914,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b01010000; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1915,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b00001010; // Expected: {'quot': 23, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1916,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 23, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1917,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b10011110; // Expected: {'quot': 1, 'rem': 71}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1918,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01100101; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1919,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1920,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 157}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1921,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1922,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011010; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011010; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1923,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1924,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b11010100; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1925,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1926,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1927,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b00011011; // Expected: {'quot': 5, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1928,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110010; Y = 8'b01010111; // Expected: {'quot': 0, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110010; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1929,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b11000011; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1930,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1931,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b10100000; // Expected: {'quot': 0, 'rem': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1932,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1933,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b00001101; // Expected: {'quot': 14, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1934,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b00100001; // Expected: {'quot': 6, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1935,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b01100101; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1936,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b00000111; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1937,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1938,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b01010100; // Expected: {'quot': 2, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1939,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1940,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1941,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000100; Y = 8'b00100000; // Expected: {'quot': 6, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000100; Y = 8'b00100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1942,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011001; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 153}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011001; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1943,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00001010; // Expected: {'quot': 12, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1944,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00111100; // Expected: {'quot': 2, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1945,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1946,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b10110001; // Expected: {'quot': 1, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1947,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b11011010; // Expected: {'quot': 0, 'rem': 189}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1948,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b01011100; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1949,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b00101110; // Expected: {'quot': 3, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1950,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b01100100; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1951,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1952,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1953,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b01010110; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1954,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b00010100; // Expected: {'quot': 10, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1955,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 223}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1956,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b00110010; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1957,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10110111; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1958,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b01101101; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b01101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1959,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b01001110; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1960,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110110; Y = 8'b00101100; // Expected: {'quot': 4, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110110; Y = 8'b00101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1961,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1962,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10000001; // Expected: {'quot': 1, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1963,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b00001111; // Expected: {'quot': 12, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1964,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b10111111; // Expected: {'quot': 0, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1965,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b00010011; // Expected: {'quot': 7, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1966,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b10010100; // Expected: {'quot': 1, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1967,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b10100001; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1968,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1969,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000010; Y = 8'b01101011; // Expected: {'quot': 1, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000010; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1970,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10000110; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1971,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b00000100; // Expected: {'quot': 37, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b00000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1972,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 37, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b10011101; // Expected: {'quot': 1, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1973,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b01000100; // Expected: {'quot': 2, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1974,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b01001100; // Expected: {'quot': 1, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1975,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b00110011; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1976,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11001010; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1977,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1978,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1979,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b00000001; // Expected: {'quot': 72, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1980,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 72, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1981,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1982,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1983,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01010101; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1984,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1985,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b10110100; // Expected: {'quot': 0, 'rem': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1986,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00001010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1987,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b01000011; // Expected: {'quot': 3, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1988,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b01101110; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1989,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1990,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b10010100; // Expected: {'quot': 1, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1991,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b00001001; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b00001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1992,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1993,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01010110; // Expected: {'quot': 2, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1994,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1995,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1996,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100010; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100010; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1997,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01010101; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1998,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b10000111; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 1999,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00000101; // Expected: {'quot': 41, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2000,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 41, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00011011; // Expected: {'quot': 8, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2001,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01100001; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2002,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b00110001; // Expected: {'quot': 3, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2003,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2004,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2005,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b00010100; // Expected: {'quot': 8, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2006,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b00111100; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2007,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2008,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b00100011; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2009,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b10000100; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b10000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2010,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b00100010; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2011,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b11011110; // Expected: {'quot': 1, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2012,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b10101010; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2013,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01111100; // Expected: {'quot': 1, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2014,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b01011000; // Expected: {'quot': 0, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b01011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2015,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010111; Y = 8'b00111101; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010111; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2016,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 138}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2017,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b11110110; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2018,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2019,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2020,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b01010011; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2021,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2022,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110111; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 55}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110111; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2023,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001110; Y = 8'b00001111; // Expected: {'quot': 0, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001110; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2024,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2025,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2026,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001001; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 73}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001001; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2027,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b00101011; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2028,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00111101; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2029,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b00010100; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b00010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2030,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10100000; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2031,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10100101; // Expected: {'quot': 1, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2032,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b10001111; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2033,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110110; Y = 8'b11101100; // Expected: {'quot': 1, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110110; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2034,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b01001111; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2035,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111010; Y = 8'b01001010; // Expected: {'quot': 0, 'rem': 58}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111010; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2036,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010001; Y = 8'b00001111; // Expected: {'quot': 9, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010001; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2037,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 137}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2038,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110101; Y = 8'b10011101; // Expected: {'quot': 0, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110101; Y = 8'b10011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2039,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b10001100; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2040,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b00111000; // Expected: {'quot': 2, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2041,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b01001101; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2042,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b01101110; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b01101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2043,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b11100011; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2044,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2045,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b00101101; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2046,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b00001111; // Expected: {'quot': 6, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2047,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 150}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2048,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b01100001; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2049,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b11011011; // Expected: {'quot': 0, 'rem': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b11011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2050,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00010010; // Expected: {'quot': 6, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2051,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2052,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b01000010; // Expected: {'quot': 3, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2053,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b10111011; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b10111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2054,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11110011; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2055,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2056,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 117}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2057,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10101111; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2058,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b00110011; // Expected: {'quot': 1, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2059,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00111000; // Expected: {'quot': 4, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2060,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2061,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01110101; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2062,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00101011; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2063,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00000101; // Expected: {'quot': 21, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2064,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 21, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10001000; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2065,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b00100010; // Expected: {'quot': 3, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2066,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b01111010; // Expected: {'quot': 0, 'rem': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2067,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010010; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010010; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2068,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b00110101; // Expected: {'quot': 4, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b00110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2069,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b01001110; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2070,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101010; Y = 8'b11010011; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101010; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2071,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b01110101; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2072,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b00100010; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2073,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b10111000; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2074,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2075,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2076,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000010; Y = 8'b10000101; // Expected: {'quot': 0, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000010; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2077,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b00110010; // Expected: {'quot': 3, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2078,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b01011011; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2079,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b10110111; // Expected: {'quot': 0, 'rem': 69}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2080,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b10011001; // Expected: {'quot': 0, 'rem': 127}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2081,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2082,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2083,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2084,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b00110100; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2085,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2086,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b01011101; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b01011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2087,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10111000; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2088,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011101; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 157}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011101; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2089,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b00010000; // Expected: {'quot': 8, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2090,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01111011; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2091,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2092,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 195}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2093,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2094,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100110; Y = 8'b11000100; // Expected: {'quot': 0, 'rem': 102}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100110; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2095,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101101; Y = 8'b10001000; // Expected: {'quot': 0, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101101; Y = 8'b10001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2096,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b10101111; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2097,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b01101011; // Expected: {'quot': 0, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2098,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111011; Y = 8'b00111100; // Expected: {'quot': 4, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111011; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2099,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2100,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00001000; // Expected: {'quot': 14, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2101,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b00000001; // Expected: {'quot': 186, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2102,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 186, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b10110101; // Expected: {'quot': 1, 'rem': 57}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2103,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2104,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2105,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10101100; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2106,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b00110100; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2107,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b00101011; // Expected: {'quot': 4, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2108,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101010; Y = 8'b10110001; // Expected: {'quot': 0, 'rem': 170}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101010; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2109,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b01100001; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2110,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b10100010; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b10100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2111,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2112,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2113,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b10011001; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2114,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b01010001; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b01010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2115,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b01100110; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2116,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 156}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2117,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2118,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01111111; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2119,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2120,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00111000; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2121,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2122,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b10101111; // Expected: {'quot': 0, 'rem': 108}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2123,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b00000101; // Expected: {'quot': 50, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2124,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 50, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b00011110; // Expected: {'quot': 5, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2125,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2126,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b00100011; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2127,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b10011011; // Expected: {'quot': 0, 'rem': 128}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2128,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b10100110; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b10100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2129,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2130,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b00001101; // Expected: {'quot': 8, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2131,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010111; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 215}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010111; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2132,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2133,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b00000011; // Expected: {'quot': 85, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b00000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2134,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 85, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b10010100; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b10010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2135,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10010000; // Expected: {'quot': 1, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2136,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2137,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b11101011; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2138,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00111110; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2139,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00100111; // Expected: {'quot': 3, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2140,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b11111010; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b11111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2141,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2142,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b10100101; // Expected: {'quot': 1, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b10100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2143,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2144,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b11010110; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2145,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b01001100; // Expected: {'quot': 3, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2146,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b10100111; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2147,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100110; Y = 8'b11001000; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100110; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2148,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2149,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b01110111; // Expected: {'quot': 1, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2150,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b10000110; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2151,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01100101; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2152,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b00001000; // Expected: {'quot': 13, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2153,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b00000001; // Expected: {'quot': 226, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2154,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2155,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2156,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b10001001; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2157,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000100; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000100; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2158,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2159,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 236}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2160,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100001; Y = 8'b01100001; // Expected: {'quot': 2, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100001; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2161,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b00101110; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2162,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2163,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111001; Y = 8'b00100011; // Expected: {'quot': 5, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111001; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2164,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b01100111; // Expected: {'quot': 2, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2165,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101100; Y = 8'b01101010; // Expected: {'quot': 1, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101100; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2166,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b01010010; // Expected: {'quot': 2, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2167,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2168,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2169,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b01011010; // Expected: {'quot': 2, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2170,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01110101; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2171,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2172,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b00101101; // Expected: {'quot': 3, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2173,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2174,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b11100011; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2175,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 132}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2176,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b01101011; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2177,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b01010001; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b01010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2178,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b00110011; // Expected: {'quot': 1, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b00110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2179,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101100; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101100; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2180,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b11000011; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2181,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2182,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b10111100; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b10111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2183,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01001000; // Expected: {'quot': 3, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2184,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b10001001; // Expected: {'quot': 0, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2185,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b00100010; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2186,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01110101; // Expected: {'quot': 1, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2187,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b00010111; // Expected: {'quot': 5, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2188,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2189,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b01010101; // Expected: {'quot': 1, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2190,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b01000111; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2191,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b00001110; // Expected: {'quot': 6, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b00001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2192,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000110; Y = 8'b00110000; // Expected: {'quot': 0, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000110; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2193,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01110100; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2194,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01000100; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2195,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000101; Y = 8'b01000000; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000101; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2196,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2197,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00010110; // Expected: {'quot': 10, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2198,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b10001010; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2199,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2200,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b10001110; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b10001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2201,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010010; Y = 8'b10110100; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010010; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2202,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b01110111; // Expected: {'quot': 1, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2203,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b00000001; // Expected: {'quot': 33, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2204,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 33, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b01001100; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2205,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000000; Y = 8'b00011010; // Expected: {'quot': 2, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000000; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2206,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 206}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2207,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 242}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2208,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2209,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00111111; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2210,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b01011001; // Expected: {'quot': 0, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2211,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01000101; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2212,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00100101; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2213,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b00010000; // Expected: {'quot': 14, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2214,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01000111; // Expected: {'quot': 2, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2215,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b01000000; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2216,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b01011100; // Expected: {'quot': 0, 'rem': 82}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2217,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b00000010; // Expected: {'quot': 78, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2218,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 78, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101100; Y = 8'b01100101; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101100; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2219,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00101110; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2220,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01001100; // Expected: {'quot': 2, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2221,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b11100100; // Expected: {'quot': 0, 'rem': 202}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b11100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2222,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b10000011; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b10000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2223,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b00100101; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b00100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2224,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b00001100; // Expected: {'quot': 19, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2225,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 19, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b10111000; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2226,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b00110100; // Expected: {'quot': 4, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2227,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b01001101; // Expected: {'quot': 2, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2228,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b10000001; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2229,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11010011; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2230,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00100100; // Expected: {'quot': 5, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2231,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b11100001; // Expected: {'quot': 0, 'rem': 152}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b11100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2232,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00101010; // Expected: {'quot': 2, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2233,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b01001101; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b01001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2234,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b01000010; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2235,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00001101; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2236,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 146}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2237,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b01010100; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2238,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00111110; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2239,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b00101011; // Expected: {'quot': 3, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2240,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b11100000; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2241,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b01010010; // Expected: {'quot': 2, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2242,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010001; Y = 8'b10101100; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010001; Y = 8'b10101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2243,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001100; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 76}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001100; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2244,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001011; Y = 8'b11000001; // Expected: {'quot': 0, 'rem': 75}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001011; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2245,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b01011001; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2246,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b00001111; // Expected: {'quot': 9, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2247,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b10010010; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2248,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 206}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2249,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111000; Y = 8'b10110011; // Expected: {'quot': 0, 'rem': 120}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111000; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2250,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2251,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b10110100; // Expected: {'quot': 0, 'rem': 70}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b10110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2252,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 124}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2253,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2254,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01100100; // Expected: {'quot': 1, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2255,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110001; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110001; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2256,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01000000; // Expected: {'quot': 2, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2257,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b01100110; // Expected: {'quot': 2, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2258,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b01000110; // Expected: {'quot': 1, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b01000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2259,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2260,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011011; Y = 8'b01000100; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011011; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2261,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b00001010; // Expected: {'quot': 23, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b00001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2262,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 23, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b10001100; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2263,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b11001010; // Expected: {'quot': 0, 'rem': 187}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b11001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2264,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b00110000; // Expected: {'quot': 1, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b00110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2265,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b10000101; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2266,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b11011000; // Expected: {'quot': 0, 'rem': 94}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2267,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101000; Y = 8'b01011001; // Expected: {'quot': 0, 'rem': 40}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101000; Y = 8'b01011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2268,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000111; Y = 8'b00000110; // Expected: {'quot': 11, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000111; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2269,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00111100; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2270,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2271,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b00011111; // Expected: {'quot': 2, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2272,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01000111; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2273,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001111; Y = 8'b10100110; // Expected: {'quot': 0, 'rem': 143}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001111; Y = 8'b10100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2274,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2275,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110100; Y = 8'b01100010; // Expected: {'quot': 1, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110100; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2276,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b01001011; // Expected: {'quot': 2, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b01001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2277,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b11111100; // Expected: {'quot': 0, 'rem': 139}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b11111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2278,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b10001010; // Expected: {'quot': 0, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b10001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2279,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b11000100; // Expected: {'quot': 0, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2280,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2281,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00100001; // Expected: {'quot': 6, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2282,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2283,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b10110001; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b10110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2284,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000100; Y = 8'b10101010; // Expected: {'quot': 0, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000100; Y = 8'b10101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2285,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00111001; // Expected: {'quot': 1, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2286,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b11000101; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2287,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111001; Y = 8'b00011111; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111001; Y = 8'b00011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2288,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 184}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2289,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b10100100; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b10100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2290,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b11011101; // Expected: {'quot': 1, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2291,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b10000001; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2292,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011101; Y = 8'b00100011; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011101; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2293,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001011; Y = 8'b00111100; // Expected: {'quot': 3, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001011; Y = 8'b00111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2294,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11100000; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2295,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b00111111; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b00111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2296,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b01011100; // Expected: {'quot': 1, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b01011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2297,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2298,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001010; Y = 8'b10011110; // Expected: {'quot': 0, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001010; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2299,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b00101110; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2300,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2301,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b10010001; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2302,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b00111101; // Expected: {'quot': 2, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b00111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2303,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100011; Y = 8'b01000011; // Expected: {'quot': 0, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100011; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2304,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2305,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b01000000; // Expected: {'quot': 3, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2306,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100010; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100010; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2307,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00000011; // Expected: {'quot': 80, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2308,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 80, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11100101; // Expected: {'quot': 0, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2309,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100101; Y = 8'b00011100; // Expected: {'quot': 8, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100101; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2310,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b01110010; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b01110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2311,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00000111; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2312,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b10110011; // Expected: {'quot': 0, 'rem': 122}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b10110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2313,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 59}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2314,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b10100001; // Expected: {'quot': 0, 'rem': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b10100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2315,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b01001010; // Expected: {'quot': 2, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2316,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2317,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b00111011; // Expected: {'quot': 2, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2318,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10010011; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2319,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b00011011; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2320,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2321,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011011; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011011; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2322,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b10010111; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2323,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b01101011; // Expected: {'quot': 0, 'rem': 105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2324,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b11011010; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b11011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2325,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b01000101; // Expected: {'quot': 1, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2326,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001110; Y = 8'b10011011; // Expected: {'quot': 1, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001110; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2327,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b01001110; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2328,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2329,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2330,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b01001010; // Expected: {'quot': 1, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b01001010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2331,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b01000001; // Expected: {'quot': 3, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2332,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b01010100; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2333,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00000110; // Expected: {'quot': 17, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2334,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b01111111; // Expected: {'quot': 1, 'rem': 68}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2335,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b01001111; // Expected: {'quot': 2, 'rem': 62}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2336,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b10010001; // Expected: {'quot': 1, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b10010001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2337,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b01110001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b01110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2338,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2339,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 126}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2340,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2341,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b11101010; // Expected: {'quot': 0, 'rem': 61}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b11101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2342,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b01100011; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2343,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b00100010; // Expected: {'quot': 7, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b00100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2344,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b00011000; // Expected: {'quot': 10, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b00011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2345,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b11101011; // Expected: {'quot': 0, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b11101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2346,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b00000010; // Expected: {'quot': 118, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b00000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2347,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 118, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b01000101; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2348,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b00011100; // Expected: {'quot': 1, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b00011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2349,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00001101; // Expected: {'quot': 8, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2350,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110101; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 181}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110101; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2351,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011011; Y = 8'b11110000; // Expected: {'quot': 0, 'rem': 219}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011011; Y = 8'b11110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2352,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110110; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 118}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110110; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2353,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000110; Y = 8'b00011011; // Expected: {'quot': 2, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000110; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2354,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2355,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100110; Y = 8'b10111001; // Expected: {'quot': 0, 'rem': 166}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100110; Y = 8'b10111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2356,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001010; Y = 8'b00010110; // Expected: {'quot': 0, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001010; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2357,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100010; Y = 8'b01101000; // Expected: {'quot': 2, 'rem': 18}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100010; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2358,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b11000100; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2359,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01000011; // Expected: {'quot': 3, 'rem': 53}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2360,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000101; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 133}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000101; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2361,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b01001011; // Expected: {'quot': 2, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b01001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2362,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b00001000; // Expected: {'quot': 6, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2363,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b00000101; // Expected: {'quot': 39, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2364,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 39, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b00010000; // Expected: {'quot': 7, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2365,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2366,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2367,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b00100111; // Expected: {'quot': 2, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b00100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2368,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b01010110; // Expected: {'quot': 2, 'rem': 66}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2369,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 131}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2370,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b10100111; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b10100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2371,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 237}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2372,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b00101011; // Expected: {'quot': 5, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2373,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b10110110; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2374,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b01110010; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b01110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2375,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2376,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00110110; // Expected: {'quot': 2, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2377,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b01011010; // Expected: {'quot': 1, 'rem': 49}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2378,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b10110010; // Expected: {'quot': 1, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2379,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100000; Y = 8'b00101111; // Expected: {'quot': 2, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100000; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2380,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b10000110; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2381,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b01111111; // Expected: {'quot': 0, 'rem': 39}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2382,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100101; Y = 8'b10100000; // Expected: {'quot': 0, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100101; Y = 8'b10100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2383,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b01100011; // Expected: {'quot': 1, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b01100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2384,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011110; Y = 8'b10101000; // Expected: {'quot': 0, 'rem': 158}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011110; Y = 8'b10101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2385,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b00011011; // Expected: {'quot': 5, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2386,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110001; Y = 8'b10111100; // Expected: {'quot': 0, 'rem': 113}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110001; Y = 8'b10111100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2387,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b11001101; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2388,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110110; Y = 8'b10111000; // Expected: {'quot': 0, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110110; Y = 8'b10111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2389,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000011; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000011; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2390,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011100; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011100; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2391,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10101101; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2392,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2393,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010011; Y = 8'b11100110; // Expected: {'quot': 0, 'rem': 147}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010011; Y = 8'b11100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2394,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101001; Y = 8'b10010111; // Expected: {'quot': 0, 'rem': 105}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101001; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2395,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b11010100; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2396,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000001; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000001; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2397,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010010; Y = 8'b00100110; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010010; Y = 8'b00100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2398,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01000001; // Expected: {'quot': 2, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2399,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01010111; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2400,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b11110001; // Expected: {'quot': 0, 'rem': 111}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b11110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2401,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b10000110; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2402,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b11010111; // Expected: {'quot': 1, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2403,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010111; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 151}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010111; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2404,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b10001100; // Expected: {'quot': 1, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2405,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b01000000; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b01000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2406,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101110; Y = 8'b11011001; // Expected: {'quot': 0, 'rem': 174}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101110; Y = 8'b11011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2407,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b01000101; // Expected: {'quot': 2, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2408,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011110; Y = 8'b01001000; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011110; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2409,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11000100; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2410,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100001; Y = 8'b00111010; // Expected: {'quot': 0, 'rem': 33}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100001; Y = 8'b00111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2411,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101001; Y = 8'b11100010; // Expected: {'quot': 0, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101001; Y = 8'b11100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2412,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111111; Y = 8'b10110101; // Expected: {'quot': 0, 'rem': 127}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111111; Y = 8'b10110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2413,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b11001111; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b11001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2414,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2415,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b10000111; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b10000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2416,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011111; Y = 8'b11001011; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011111; Y = 8'b11001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2417,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011110; Y = 8'b00101111; // Expected: {'quot': 0, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011110; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2418,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b10001100; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b10001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2419,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2420,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b10011100; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b10011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2421,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011111; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011111; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2422,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b01001111; // Expected: {'quot': 2, 'rem': 10}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2423,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b00100000; // Expected: {'quot': 6, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b00100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2424,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101111; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101111; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2425,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101101; Y = 8'b01101011; // Expected: {'quot': 1, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101101; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2426,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2427,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b00100000; // Expected: {'quot': 7, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b00100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2428,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101011; Y = 8'b11000001; // Expected: {'quot': 1, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101011; Y = 8'b11000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2429,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011100; Y = 8'b11110110; // Expected: {'quot': 0, 'rem': 220}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011100; Y = 8'b11110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2430,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 244}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2431,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000000; Y = 8'b11011111; // Expected: {'quot': 0, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000000; Y = 8'b11011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2432,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b00110100; // Expected: {'quot': 4, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b00110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2433,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b11110111; // Expected: {'quot': 0, 'rem': 212}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b11110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2434,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011000; Y = 8'b11001000; // Expected: {'quot': 0, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011000; Y = 8'b11001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2435,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00111011; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2436,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b01110110; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2437,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b00100011; // Expected: {'quot': 3, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b00100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2438,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001101; Y = 8'b01100111; // Expected: {'quot': 0, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001101; Y = 8'b01100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2439,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010101; Y = 8'b01111001; // Expected: {'quot': 0, 'rem': 85}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010101; Y = 8'b01111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2440,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100000; Y = 8'b11000000; // Expected: {'quot': 1, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100000; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2441,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101000; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 168}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101000; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2442,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2443,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b11101111; // Expected: {'quot': 0, 'rem': 162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2444,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01110011; // Expected: {'quot': 1, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2445,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001011; Y = 8'b01101011; // Expected: {'quot': 0, 'rem': 11}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001011; Y = 8'b01101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2446,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b11001110; // Expected: {'quot': 0, 'rem': 190}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b11001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2447,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b11010101; // Expected: {'quot': 0, 'rem': 84}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b11010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2448,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101111; Y = 8'b10011110; // Expected: {'quot': 1, 'rem': 81}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101111; Y = 8'b10011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2449,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b00010011; // Expected: {'quot': 2, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b00010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2450,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b00110001; // Expected: {'quot': 1, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2451,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111000; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111000; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2452,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b01011011; // Expected: {'quot': 2, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b01011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2453,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b01111000; // Expected: {'quot': 1, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2454,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b11010110; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b11010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2455,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b01100010; // Expected: {'quot': 0, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b01100010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2456,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110001; Y = 8'b10010010; // Expected: {'quot': 1, 'rem': 95}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110001; Y = 8'b10010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2457,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2458,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111110; Y = 8'b10011001; // Expected: {'quot': 1, 'rem': 37}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111110; Y = 8'b10011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2459,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011010; Y = 8'b01000011; // Expected: {'quot': 3, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011010; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2460,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 178}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2461,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011001; Y = 8'b11101110; // Expected: {'quot': 0, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011001; Y = 8'b11101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2462,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b01001111; // Expected: {'quot': 2, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b01001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2463,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000000; Y = 8'b00010111; // Expected: {'quot': 5, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000000; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2464,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100000; Y = 8'b10000110; // Expected: {'quot': 1, 'rem': 26}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100000; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2465,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b11011000; // Expected: {'quot': 1, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2466,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b11101000; // Expected: {'quot': 0, 'rem': 149}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b11101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2467,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101111; Y = 8'b01000001; // Expected: {'quot': 2, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101111; Y = 8'b01000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2468,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01000011; // Expected: {'quot': 3, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2469,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101100; Y = 8'b11001100; // Expected: {'quot': 1, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101100; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2470,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b10011000; // Expected: {'quot': 1, 'rem': 98}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b10011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2471,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b10000010; // Expected: {'quot': 1, 'rem': 77}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2472,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b01100110; // Expected: {'quot': 1, 'rem': 74}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b01100110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2473,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11001101; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2474,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001101; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 205}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001101; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2475,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b00101110; // Expected: {'quot': 2, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b00101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2476,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101101; Y = 8'b00100001; // Expected: {'quot': 7, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101101; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2477,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110011; Y = 8'b11101111; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110011; Y = 8'b11101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2478,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2479,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b00110010; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b00110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2480,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111101; Y = 8'b00110001; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111101; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2481,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100011; Y = 8'b01010010; // Expected: {'quot': 2, 'rem': 63}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100011; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2482,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100010; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 162}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100010; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2483,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100110; Y = 8'b00000001; // Expected: {'quot': 38, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100110; Y = 8'b00000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2484,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 38, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010110; Y = 8'b01000101; // Expected: {'quot': 2, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010110; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2485,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001001; Y = 8'b00100001; // Expected: {'quot': 4, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001001; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2486,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110111; Y = 8'b10010110; // Expected: {'quot': 1, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110111; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2487,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 140}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2488,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10010000; // Expected: {'quot': 1, 'rem': 44}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2489,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101110; Y = 8'b11111000; // Expected: {'quot': 0, 'rem': 110}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101110; Y = 8'b11111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2490,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b11000110; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b11000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2491,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b00011001; // Expected: {'quot': 7, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b00011001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2492,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b01101000; // Expected: {'quot': 2, 'rem': 47}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2493,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011110; Y = 8'b00011011; // Expected: {'quot': 8, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011110; Y = 8'b00011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2494,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011010; Y = 8'b11110100; // Expected: {'quot': 0, 'rem': 154}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011010; Y = 8'b11110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2495,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010001; Y = 8'b00101111; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010001; Y = 8'b00101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2496,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100111; Y = 8'b00011101; // Expected: {'quot': 7, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100111; Y = 8'b00011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2497,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111111; Y = 8'b01110100; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111111; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2498,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b01001011; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b01001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2499,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111001; Y = 8'b10001011; // Expected: {'quot': 0, 'rem': 121}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111001; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2500,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b10101110; // Expected: {'quot': 1, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2501,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011001; Y = 8'b00010110; // Expected: {'quot': 9, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011001; Y = 8'b00010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2502,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000111; Y = 8'b10010101; // Expected: {'quot': 0, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000111; Y = 8'b10010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2503,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111010; Y = 8'b11110011; // Expected: {'quot': 1, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111010; Y = 8'b11110011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2504,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010100; Y = 8'b00101001; // Expected: {'quot': 3, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010100; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2505,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01101000; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2506,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b00111000; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b00111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2507,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101010; Y = 8'b11111110; // Expected: {'quot': 0, 'rem': 42}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101010; Y = 8'b11111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2508,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010111; Y = 8'b01011010; // Expected: {'quot': 0, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010111; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2509,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110010; Y = 8'b01010101; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110010; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2510,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001110; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 142}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001110; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2511,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b11111111; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b11111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2512,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b01000010; // Expected: {'quot': 1, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2513,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00000101; // Expected: {'quot': 11, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2514,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111011; Y = 8'b00010111; // Expected: {'quot': 5, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111011; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2515,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b00111001; // Expected: {'quot': 3, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2516,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b10010111; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b10010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2517,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b11101001; // Expected: {'quot': 0, 'rem': 228}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b11101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2518,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100100; Y = 8'b01110100; // Expected: {'quot': 0, 'rem': 36}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100100; Y = 8'b01110100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2519,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010000; Y = 8'b00010000; // Expected: {'quot': 5, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010000; Y = 8'b00010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2520,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110100; Y = 8'b01011111; // Expected: {'quot': 2, 'rem': 54}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110100; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2521,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00010101; // Expected: {'quot': 8, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2522,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101000; Y = 8'b01000101; // Expected: {'quot': 3, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101000; Y = 8'b01000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2523,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b01111110; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b01111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2524,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b11001001; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2525,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b01110111; // Expected: {'quot': 1, 'rem': 64}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2526,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111011; Y = 8'b00001111; // Expected: {'quot': 3, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111011; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2527,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111111; Y = 8'b00100001; // Expected: {'quot': 1, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111111; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2528,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b01000111; // Expected: {'quot': 2, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2529,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000111; Y = 8'b01010101; // Expected: {'quot': 2, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000111; Y = 8'b01010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2530,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110000; Y = 8'b01010100; // Expected: {'quot': 1, 'rem': 28}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110000; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2531,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110101; Y = 8'b00101001; // Expected: {'quot': 2, 'rem': 35}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110101; Y = 8'b00101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2532,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011000; Y = 8'b00000111; // Expected: {'quot': 21, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011000; Y = 8'b00000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2533,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 21, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101001; Y = 8'b01010011; // Expected: {'quot': 2, 'rem': 3}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101001; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2534,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00111001; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2535,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110011; Y = 8'b10111101; // Expected: {'quot': 0, 'rem': 179}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110011; Y = 8'b10111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2536,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b00001100; // Expected: {'quot': 14, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2537,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b00010111; // Expected: {'quot': 7, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2538,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 7, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b11110010; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b11110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2539,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111000; Y = 8'b00001111; // Expected: {'quot': 12, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111000; Y = 8'b00001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2540,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 12, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2541,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011111; Y = 8'b01101001; // Expected: {'quot': 0, 'rem': 31}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011111; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2542,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 80}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2543,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010101; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 149}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010101; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2544,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010011; Y = 8'b10110110; // Expected: {'quot': 1, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010011; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2545,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110100; Y = 8'b00001000; // Expected: {'quot': 22, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110100; Y = 8'b00001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2546,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 22, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b00100100; // Expected: {'quot': 6, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b00100100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2547,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111011; Y = 8'b10101110; // Expected: {'quot': 1, 'rem': 13}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111011; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2548,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001000; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001000; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2549,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b11010010; // Expected: {'quot': 0, 'rem': 141}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b11010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2550,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111110; Y = 8'b01110101; // Expected: {'quot': 1, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111110; Y = 8'b01110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2551,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010100; Y = 8'b10111111; // Expected: {'quot': 1, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010100; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2552,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110000; Y = 8'b01101000; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110000; Y = 8'b01101000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2553,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000100; Y = 8'b01111111; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000100; Y = 8'b01111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2554,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000101; Y = 8'b01101010; // Expected: {'quot': 1, 'rem': 91}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000101; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2555,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010110; Y = 8'b00000110; // Expected: {'quot': 35, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010110; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2556,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 35, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011011; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011011; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2557,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110100; Y = 8'b11011100; // Expected: {'quot': 0, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110100; Y = 8'b11011100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2558,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001100; Y = 8'b11100011; // Expected: {'quot': 0, 'rem': 204}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001100; Y = 8'b11100011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2559,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b11011101; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b11011101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2560,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b00010111; // Expected: {'quot': 6, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b00010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2561,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111001; Y = 8'b00011010; // Expected: {'quot': 9, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111001; Y = 8'b00011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2562,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111101; Y = 8'b10010011; // Expected: {'quot': 1, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111101; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2563,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b00000110; // Expected: {'quot': 17, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b00000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2564,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 17, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011010; Y = 8'b11101100; // Expected: {'quot': 0, 'rem': 90}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011010; Y = 8'b11101100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2565,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110001; Y = 8'b10001011; // Expected: {'quot': 1, 'rem': 38}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110001; Y = 8'b10001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2566,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010001; Y = 8'b11001100; // Expected: {'quot': 0, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010001; Y = 8'b11001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2567,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b00111011; // Expected: {'quot': 1, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2568,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110011; Y = 8'b10111010; // Expected: {'quot': 0, 'rem': 51}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110011; Y = 8'b10111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2569,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001110; Y = 8'b01011010; // Expected: {'quot': 0, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001110; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2570,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100100; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 100}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100100; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2571,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010110; Y = 8'b00110001; // Expected: {'quot': 0, 'rem': 22}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010110; Y = 8'b00110001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2572,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010000; Y = 8'b11010011; // Expected: {'quot': 0, 'rem': 16}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010000; Y = 8'b11010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2573,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001100; Y = 8'b01011111; // Expected: {'quot': 0, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001100; Y = 8'b01011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2574,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111010; Y = 8'b00111001; // Expected: {'quot': 2, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111010; Y = 8'b00111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2575,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000110; Y = 8'b11001001; // Expected: {'quot': 0, 'rem': 198}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000110; Y = 8'b11001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2576,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010011; Y = 8'b01111000; // Expected: {'quot': 0, 'rem': 83}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010011; Y = 8'b01111000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2577,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101000; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 104}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101000; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2578,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111000; Y = 8'b10011011; // Expected: {'quot': 1, 'rem': 93}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111000; Y = 8'b10011011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2579,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001100; Y = 8'b01011010; // Expected: {'quot': 1, 'rem': 50}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001100; Y = 8'b01011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2580,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10101011; Y = 8'b11010000; // Expected: {'quot': 0, 'rem': 171}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10101011; Y = 8'b11010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2581,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000001; Y = 8'b11000101; // Expected: {'quot': 0, 'rem': 129}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000001; Y = 8'b11000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2582,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10011010; // Expected: {'quot': 1, 'rem': 34}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10011010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2583,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111111; Y = 8'b10111111; // Expected: {'quot': 1, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111111; Y = 8'b10111111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2584,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10110010; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10110010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2585,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110000; Y = 8'b11011000; // Expected: {'quot': 1, 'rem': 24}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110000; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2586,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001111; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001111; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2587,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001101; Y = 8'b10001001; // Expected: {'quot': 1, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001101; Y = 8'b10001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2588,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000010; Y = 8'b01010000; // Expected: {'quot': 0, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000010; Y = 8'b01010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2589,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111100; Y = 8'b10001111; // Expected: {'quot': 1, 'rem': 45}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111100; Y = 8'b10001111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2590,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 99}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2591,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101010; Y = 8'b01110111; // Expected: {'quot': 0, 'rem': 106}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101010; Y = 8'b01110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2592,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b01000010; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b01000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2593,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100000; Y = 8'b01101010; // Expected: {'quot': 0, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100000; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2594,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b01111010; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b01111010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2595,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111101; Y = 8'b10101111; // Expected: {'quot': 1, 'rem': 14}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111101; Y = 8'b10101111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2596,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b11000011; // Expected: {'quot': 0, 'rem': 89}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b11000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2597,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111100; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111100; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2598,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001000; Y = 8'b11000010; // Expected: {'quot': 0, 'rem': 136}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001000; Y = 8'b11000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2599,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011000; Y = 8'b11011000; // Expected: {'quot': 0, 'rem': 88}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011000; Y = 8'b11011000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2600,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001111; Y = 8'b00111011; // Expected: {'quot': 3, 'rem': 30}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001111; Y = 8'b00111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2601,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010011; Y = 8'b10101001; // Expected: {'quot': 0, 'rem': 19}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010011; Y = 8'b10101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2602,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100101; Y = 8'b11111001; // Expected: {'quot': 0, 'rem': 101}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100101; Y = 8'b11111001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2603,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b01000100; // Expected: {'quot': 1, 'rem': 56}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b01000100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2604,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11100100; Y = 8'b01000011; // Expected: {'quot': 3, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11100100; Y = 8'b01000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2605,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b01010110; // Expected: {'quot': 1, 'rem': 17}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b01010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2606,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000111; Y = 8'b10111110; // Expected: {'quot': 0, 'rem': 135}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000111; Y = 8'b10111110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2607,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111100; Y = 8'b00001101; // Expected: {'quot': 9, 'rem': 7}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111100; Y = 8'b00001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2608,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110010; Y = 8'b01010010; // Expected: {'quot': 2, 'rem': 78}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110010; Y = 8'b01010010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2609,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101110; Y = 8'b11111011; // Expected: {'quot': 0, 'rem': 238}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101110; Y = 8'b11111011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2610,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11111110; Y = 8'b01100101; // Expected: {'quot': 2, 'rem': 52}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11111110; Y = 8'b01100101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2611,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01001111; Y = 8'b11100111; // Expected: {'quot': 0, 'rem': 79}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01001111; Y = 8'b11100111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2612,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010110; Y = 8'b11101101; // Expected: {'quot': 0, 'rem': 86}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010110; Y = 8'b11101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2613,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001011; Y = 8'b01001000; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001011; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2614,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00011101; Y = 8'b01100000; // Expected: {'quot': 0, 'rem': 29}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00011101; Y = 8'b01100000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2615,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101011; Y = 8'b01110000; // Expected: {'quot': 0, 'rem': 43}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101011; Y = 8'b01110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2616,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10111010; Y = 8'b11011110; // Expected: {'quot': 0, 'rem': 186}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10111010; Y = 8'b11011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2617,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000001; Y = 8'b01010011; // Expected: {'quot': 2, 'rem': 27}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000001; Y = 8'b01010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2618,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b01100001; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b01100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2619,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01000001; Y = 8'b10000010; // Expected: {'quot': 0, 'rem': 65}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01000001; Y = 8'b10000010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2620,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101011; Y = 8'b10011111; // Expected: {'quot': 0, 'rem': 107}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101011; Y = 8'b10011111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2621,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00101110; Y = 8'b10010110; // Expected: {'quot': 0, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00101110; Y = 8'b10010110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2622,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000000; Y = 8'b11010100; // Expected: {'quot': 0, 'rem': 192}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000000; Y = 8'b11010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2623,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010000; Y = 8'b10101110; // Expected: {'quot': 0, 'rem': 144}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010000; Y = 8'b10101110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2624,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10001010; Y = 8'b01101010; // Expected: {'quot': 1, 'rem': 32}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10001010; Y = 8'b01101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2625,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11101001; Y = 8'b10101101; // Expected: {'quot': 1, 'rem': 60}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11101001; Y = 8'b10101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2626,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100111; Y = 8'b10110110; // Expected: {'quot': 0, 'rem': 167}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100111; Y = 8'b10110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2627,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11000011; Y = 8'b10010101; // Expected: {'quot': 1, 'rem': 46}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11000011; Y = 8'b10010101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2628,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001010; Y = 8'b00100001; // Expected: {'quot': 6, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001010; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2629,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01010100; Y = 8'b01001000; // Expected: {'quot': 1, 'rem': 12}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01010100; Y = 8'b01001000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2630,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01110111; Y = 8'b11111101; // Expected: {'quot': 0, 'rem': 119}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01110111; Y = 8'b11111101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2631,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00100111; Y = 8'b00001011; // Expected: {'quot': 3, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00100111; Y = 8'b00001011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2632,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10010010; Y = 8'b01000111; // Expected: {'quot': 2, 'rem': 4}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10010010; Y = 8'b01000111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2633,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100100; Y = 8'b10110111; // Expected: {'quot': 0, 'rem': 164}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100100; Y = 8'b10110111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2634,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100101; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 165}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100101; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2635,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000110; Y = 8'b10000001; // Expected: {'quot': 1, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000110; Y = 8'b10000001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2636,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00000101; Y = 8'b10010011; // Expected: {'quot': 0, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00000101; Y = 8'b10010011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2637,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100011; Y = 8'b01010100; // Expected: {'quot': 1, 'rem': 15}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100011; Y = 8'b01010100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2638,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001000; Y = 8'b10010000; // Expected: {'quot': 0, 'rem': 8}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001000; Y = 8'b10010000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2639,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10000011; Y = 8'b00101010; // Expected: {'quot': 3, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10000011; Y = 8'b00101010; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2640,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00110000; Y = 8'b01001001; // Expected: {'quot': 0, 'rem': 48}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00110000; Y = 8'b01001001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2641,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10100011; Y = 8'b00000011; // Expected: {'quot': 54, 'rem': 1}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10100011; Y = 8'b00000011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2642,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 54, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11010101; Y = 8'b10001101; // Expected: {'quot': 1, 'rem': 72}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11010101; Y = 8'b10001101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2643,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01011001; Y = 8'b00100001; // Expected: {'quot': 2, 'rem': 23}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01011001; Y = 8'b00100001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2644,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010101; Y = 8'b11110101; // Expected: {'quot': 0, 'rem': 21}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010101; Y = 8'b11110101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2645,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011101; Y = 8'b10000110; // Expected: {'quot': 1, 'rem': 87}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011101; Y = 8'b10000110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2646,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11011000; Y = 8'b01101001; // Expected: {'quot': 2, 'rem': 6}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11011000; Y = 8'b01101001; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2647,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01111101; Y = 8'b10000000; // Expected: {'quot': 0, 'rem': 125}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01111101; Y = 8'b10000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2648,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11001000; Y = 8'b10000101; // Expected: {'quot': 1, 'rem': 67}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11001000; Y = 8'b10000101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2649,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011111; Y = 8'b01110110; // Expected: {'quot': 1, 'rem': 41}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011111; Y = 8'b01110110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2650,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 1, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100001; Y = 8'b11000000; // Expected: {'quot': 0, 'rem': 97}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100001; Y = 8'b11000000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2651,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01101111; Y = 8'b00101011; // Expected: {'quot': 2, 'rem': 25}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01101111; Y = 8'b00101011; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2652,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b01100111; Y = 8'b10110000; // Expected: {'quot': 0, 'rem': 103}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b01100111; Y = 8'b10110000; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2653,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00111110; Y = 8'b00001100; // Expected: {'quot': 5, 'rem': 2}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00111110; Y = 8'b00001100; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2654,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10011100; Y = 8'b01001110; // Expected: {'quot': 2, 'rem': 0}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10011100; Y = 8'b01001110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2655,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b10110111; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 183}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b10110111; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2656,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00001001; Y = 8'b11010111; // Expected: {'quot': 0, 'rem': 9}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00001001; Y = 8'b11010111; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2657,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b00010100; Y = 8'b00101101; // Expected: {'quot': 0, 'rem': 20}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b00010100; Y = 8'b00101101; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2658,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 0, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 X = 8'b11110101; Y = 8'b00011110; // Expected: {'quot': 8, 'rem': 5}
        
        start = 1'b1;
        #10 start = 1'b0;
        
        
        wait(valid);
        
        
        $display("Test %0d: Inputs: X = 8'b11110101; Y = 8'b00011110; | Outputs: quot=%b, rem=%b, valid=%b | Expected: quot=%d, rem=%d",
                 2659,
                 
                 quot, 
                 
                 rem, 
                 
                 valid
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule