
`timescale 1ns / 1ps

module tb_N8_carry_save_adder_l2;

    // Parameters
    
    parameter N = 8;
    
     
    // Inputs
    
    reg  [7:0] a;
    
    reg  [7:0] b;
    
    reg  [7:0] c;
    
    
    // Outputs
    
    wire  [7:0] sum;
    
    wire  [7:0] carry;
    
    
    // Instantiate the Unit Under Test (UUT)
    carry_save_adder_l2  #( N ) uut (
        
        .a(a),
        
        .b(b),
        
        .c(c),
        
        
        .sum(sum),
        
        .carry(carry)
        
    );
    
    initial begin
        // Initialize Inputs
        
        a = 0;
        
        b = 0;
        
        c = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        a = 8'b10101001; b = 8'b01111000; c = 8'b00011011; // Expected: {'sum': 202, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01111000; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 0,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b01101010; c = 8'b10110101; // Expected: {'sum': 81, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b01101010; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00101100; c = 8'b01101111; // Expected: {'sum': 3, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00101100; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00100011; c = 8'b00101010; // Expected: {'sum': 231, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00100011; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11110000; c = 8'b01101011; // Expected: {'sum': 73, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11110000; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 4,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00010001; c = 8'b01111011; // Expected: {'sum': 31, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00010001; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 5,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00110101; c = 8'b11100110; // Expected: {'sum': 215, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00110101; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 6,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11010101; c = 8'b01000011; // Expected: {'sum': 72, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11010101; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 7,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01101111; c = 8'b01011110; // Expected: {'sum': 228, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01101111; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 8,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b11000000; c = 8'b01111100; // Expected: {'sum': 161, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b11000000; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 9,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11000110; c = 8'b10111001; // Expected: {'sum': 134, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11000110; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 10,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b01111000; c = 8'b10111110; // Expected: {'sum': 33, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b01111000; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 11,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10101011; c = 8'b11000011; // Expected: {'sum': 123, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10101011; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 12,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b10010101; c = 8'b10000001; // Expected: {'sum': 97, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b10010101; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 13,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01000101; c = 8'b01001001; // Expected: {'sum': 122, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01000101; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 14,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00110101; c = 8'b10110101; // Expected: {'sum': 174, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00110101; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 15,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00011111; c = 8'b00010011; // Expected: {'sum': 113, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00011111; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 16,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11010110; c = 8'b10110010; // Expected: {'sum': 53, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11010110; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 17,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01000101; c = 8'b11100000; // Expected: {'sum': 159, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01000101; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 18,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11011011; c = 8'b01100111; // Expected: {'sum': 158, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11011011; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 19,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10011110; c = 8'b10010111; // Expected: {'sum': 191, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10011110; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 20,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01011100; c = 8'b00111110; // Expected: {'sum': 10, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01011100; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 21,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01110011; c = 8'b01011011; // Expected: {'sum': 52, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01110011; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 22,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00001100; c = 8'b00010111; // Expected: {'sum': 45, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00001100; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 23,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10001001; c = 8'b10011101; // Expected: {'sum': 169, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10001001; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 24,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10100000; c = 8'b00100001; // Expected: {'sum': 75, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10100000; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 25,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11000000; c = 8'b10110000; // Expected: {'sum': 136, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11000000; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 26,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00000001; c = 8'b11011000; // Expected: {'sum': 72, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00000001; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 27,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10011010; c = 8'b11101101; // Expected: {'sum': 173, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10011010; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 28,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01001110; c = 8'b01001101; // Expected: {'sum': 144, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01001110; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 29,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01001111; c = 8'b00001100; // Expected: {'sum': 61, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01001111; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 30,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00111010; c = 8'b11110100; // Expected: {'sum': 10, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00111010; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 31,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b10000111; c = 8'b10110011; // Expected: {'sum': 124, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b10000111; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 32,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10011101; c = 8'b01010100; // Expected: {'sum': 255, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10011101; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 33,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00100101; c = 8'b10000110; // Expected: {'sum': 231, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00100101; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 34,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b11111010; c = 8'b11010010; // Expected: {'sum': 56, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b11111010; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 35,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10100011; c = 8'b01111100; // Expected: {'sum': 81, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10100011; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 36,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00001000; c = 8'b10101010; // Expected: {'sum': 197, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00001000; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 37,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00001010; c = 8'b01000111; // Expected: {'sum': 183, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00001010; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 38,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b10110110; c = 8'b10101001; // Expected: {'sum': 42, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b10110110; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 39,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01111110; c = 8'b00110110; // Expected: {'sum': 73, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01111110; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 40,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11011100; c = 8'b01010101; // Expected: {'sum': 38, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11011100; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 41,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00001101; c = 8'b11110100; // Expected: {'sum': 111, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00001101; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 42,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00101100; c = 8'b11011111; // Expected: {'sum': 237, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00101100; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 43,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00011011; c = 8'b10001111; // Expected: {'sum': 118, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00011011; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 44,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10010001; c = 8'b01011110; // Expected: {'sum': 112, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10010001; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 45,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10110000; c = 8'b00000010; // Expected: {'sum': 90, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10110000; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 46,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10110010; c = 8'b00001011; // Expected: {'sum': 179, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10110010; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 47,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10100100; c = 8'b01110000; // Expected: {'sum': 69, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10100100; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 48,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b00011111; c = 8'b11101100; // Expected: {'sum': 139, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b00011111; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 49,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01000010; c = 8'b00100010; // Expected: {'sum': 146, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01000010; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 50,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10100001; c = 8'b01111000; // Expected: {'sum': 214, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10100001; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 51,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00010111; c = 8'b01011100; // Expected: {'sum': 176, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00010111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 52,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b11000001; c = 8'b01011100; // Expected: {'sum': 197, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b11000001; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 53,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01100100; c = 8'b11000000; // Expected: {'sum': 164, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01100100; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 54,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11111110; c = 8'b11000001; // Expected: {'sum': 66, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11111110; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 55,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b00010010; c = 8'b01101001; // Expected: {'sum': 254, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b00010010; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 56,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11111010; c = 8'b00101100; // Expected: {'sum': 180, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11111010; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 57,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01100101; c = 8'b10100110; // Expected: {'sum': 51, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01100101; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 58,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11100100; c = 8'b10011011; // Expected: {'sum': 205, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11100100; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 59,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10000001; c = 8'b10100010; // Expected: {'sum': 78, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10000001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 60,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00101110; c = 8'b10111010; // Expected: {'sum': 237, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00101110; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 61,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11100011; c = 8'b10000011; // Expected: {'sum': 73, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11100011; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 62,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b01000100; c = 8'b00110011; // Expected: {'sum': 98, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b01000100; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 63,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10100010; c = 8'b11110100; // Expected: {'sum': 69, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10100010; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 64,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00001010; c = 8'b01100000; // Expected: {'sum': 115, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00001010; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 65,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b00110101; c = 8'b11100100; // Expected: {'sum': 119, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b00110101; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 66,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b01101111; c = 8'b10101111; // Expected: {'sum': 103, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b01101111; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 67,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00000010; c = 8'b11110011; // Expected: {'sum': 15, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00000010; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 68,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01110001; c = 8'b01010000; // Expected: {'sum': 21, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01110001; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 69,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10000010; c = 8'b01011010; // Expected: {'sum': 49, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10000010; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 70,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01011010; c = 8'b11100011; // Expected: {'sum': 76, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01011010; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 71,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10001011; c = 8'b01111000; // Expected: {'sum': 98, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10001011; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 72,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00010001; c = 8'b01100010; // Expected: {'sum': 152, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00010001; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 73,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11101001; c = 8'b01000100; // Expected: {'sum': 86, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11101001; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 74,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00111000; c = 8'b01000101; // Expected: {'sum': 10, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00111000; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 75,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00111101; c = 8'b10001101; // Expected: {'sum': 153, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00111101; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 76,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11000100; c = 8'b11100111; // Expected: {'sum': 128, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11000100; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 77,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10110010; c = 8'b00100010; // Expected: {'sum': 51, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10110010; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 78,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00111001; c = 8'b01111101; // Expected: {'sum': 138, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00111001; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 79,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01101000; c = 8'b01101001; // Expected: {'sum': 151, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01101000; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 80,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10111011; c = 8'b00111011; // Expected: {'sum': 244, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10111011; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 81,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01100001; c = 8'b00110101; // Expected: {'sum': 112, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01100001; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 82,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00101110; c = 8'b01001111; // Expected: {'sum': 240, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00101110; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 83,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10101010; c = 8'b10001110; // Expected: {'sum': 176, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10101010; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 84,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01011111; c = 8'b01011101; // Expected: {'sum': 236, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01011111; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 85,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11000010; c = 8'b01110111; // Expected: {'sum': 209, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11000010; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 86,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b11111000; c = 8'b01010111; // Expected: {'sum': 14, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b11111000; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 87,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00111001; c = 8'b00100101; // Expected: {'sum': 240, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00111001; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 88,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11110110; c = 8'b00000001; // Expected: {'sum': 2, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11110110; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 89,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10100101; c = 8'b11001110; // Expected: {'sum': 233, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10100101; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 90,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00100100; c = 8'b11100111; // Expected: {'sum': 108, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00100100; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 91,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00101100; c = 8'b00111100; // Expected: {'sum': 208, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00101100; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 92,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b00011110; c = 8'b10011101; // Expected: {'sum': 82, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b00011110; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 93,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b01011100; c = 8'b01001100; // Expected: {'sum': 146, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b01011100; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 94,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10100010; c = 8'b00111001; // Expected: {'sum': 75, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10100010; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 95,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b11010000; c = 8'b11010000; // Expected: {'sum': 156, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b11010000; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 96,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b10111010; c = 8'b00011111; // Expected: {'sum': 88, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b10111010; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 97,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01110111; c = 8'b00010011; // Expected: {'sum': 220, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01110111; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 98,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01001101; c = 8'b00000011; // Expected: {'sum': 132, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01001101; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 99,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10110101; c = 8'b01100000; // Expected: {'sum': 14, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10110101; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10111000; c = 8'b00100110; // Expected: {'sum': 4, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10111000; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01011110; c = 8'b11101111; // Expected: {'sum': 85, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01011110; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b11111000; c = 8'b01101010; // Expected: {'sum': 245, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b11111000; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11000010; c = 8'b00010010; // Expected: {'sum': 226, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11000010; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11010011; c = 8'b10111110; // Expected: {'sum': 233, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11010011; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b11000100; c = 8'b01000101; // Expected: {'sum': 188, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b11000100; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10001000; c = 8'b11001010; // Expected: {'sum': 66, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10001000; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10011100; c = 8'b01010110; // Expected: {'sum': 112, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10011100; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11101100; c = 8'b01010001; // Expected: {'sum': 171, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11101100; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11101101; c = 8'b10010001; // Expected: {'sum': 235, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11101101; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00010100; c = 8'b10110100; // Expected: {'sum': 59, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00010100; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10111001; c = 8'b11100110; // Expected: {'sum': 143, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10111001; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11101110; c = 8'b01011011; // Expected: {'sum': 102, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11101110; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b01111010; c = 8'b10100101; // Expected: {'sum': 211, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b01111010; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b01000001; c = 8'b11110001; // Expected: {'sum': 185, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b01000001; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b01111101; c = 8'b00010100; // Expected: {'sum': 243, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b01111101; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10101010; c = 8'b10110001; // Expected: {'sum': 11, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10101010; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00001101; c = 8'b00101000; // Expected: {'sum': 128, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00001101; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10011011; c = 8'b01001101; // Expected: {'sum': 5, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10011011; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10111110; c = 8'b00001000; // Expected: {'sum': 11, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10111110; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01110111; c = 8'b01011100; // Expected: {'sum': 12, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01110111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00111100; c = 8'b01111001; // Expected: {'sum': 190, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00111100; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b10000100; c = 8'b00111110; // Expected: {'sum': 243, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b10000100; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10011000; c = 8'b00101111; // Expected: {'sum': 52, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10011000; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01100111; c = 8'b11111101; // Expected: {'sum': 19, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01100111; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11011100; c = 8'b11110001; // Expected: {'sum': 71, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11011100; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11110101; c = 8'b00110111; // Expected: {'sum': 87, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11110101; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b10011101; c = 8'b11000110; // Expected: {'sum': 205, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b10011101; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01011000; c = 8'b01001111; // Expected: {'sum': 158, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01011000; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11000111; c = 8'b00010000; // Expected: {'sum': 74, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11000111; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11110011; c = 8'b00101010; // Expected: {'sum': 85, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11110011; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11111011; c = 8'b10001101; // Expected: {'sum': 196, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11111011; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b11100100; c = 8'b00011101; // Expected: {'sum': 21, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b11100100; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11100011; c = 8'b00010011; // Expected: {'sum': 190, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11100011; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11111111; c = 8'b10010000; // Expected: {'sum': 24, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11111111; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b11000110; c = 8'b10101111; // Expected: {'sum': 230, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b11000110; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b10011111; c = 8'b11101100; // Expected: {'sum': 66, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b10011111; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01010011; c = 8'b00000011; // Expected: {'sum': 195, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01010011; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01100011; c = 8'b00100000; // Expected: {'sum': 117, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01100011; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10000111; c = 8'b01101100; // Expected: {'sum': 250, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10000111; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b11101010; c = 8'b10101010; // Expected: {'sum': 16, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b11101010; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01011011; c = 8'b11011110; // Expected: {'sum': 115, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01011011; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01101110; c = 8'b00011001; // Expected: {'sum': 52, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01101110; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10000011; c = 8'b11000011; // Expected: {'sum': 185, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10000011; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10010010; c = 8'b11110111; // Expected: {'sum': 221, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10010010; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11111000; c = 8'b01011100; // Expected: {'sum': 63, 'carry': 216}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11111000; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00001100; c = 8'b00111010; // Expected: {'sum': 123, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00001100; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01011001; c = 8'b00101101; // Expected: {'sum': 12, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01011001; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01111101; c = 8'b10100011; // Expected: {'sum': 6, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01111101; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10111001; c = 8'b11110000; // Expected: {'sum': 127, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10111001; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11000100; c = 8'b10110101; // Expected: {'sum': 125, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11000100; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01000110; c = 8'b01101100; // Expected: {'sum': 204, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01000110; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11111110; c = 8'b10011000; // Expected: {'sum': 130, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11111110; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10000101; c = 8'b11011101; // Expected: {'sum': 252, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10000101; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10010110; c = 8'b01100001; // Expected: {'sum': 3, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10010110; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00110001; c = 8'b00111100; // Expected: {'sum': 185, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00110001; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11001111; c = 8'b10000100; // Expected: {'sum': 227, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11001111; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00000010; c = 8'b11100111; // Expected: {'sum': 146, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00000010; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11000110; c = 8'b00001011; // Expected: {'sum': 84, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11000110; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01100110; c = 8'b10100111; // Expected: {'sum': 78, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01100110; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00010100; c = 8'b00110111; // Expected: {'sum': 217, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00010100; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b11001100; c = 8'b01101100; // Expected: {'sum': 233, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b11001100; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10011101; c = 8'b00011110; // Expected: {'sum': 173, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10011101; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b01010000; c = 8'b00010000; // Expected: {'sum': 66, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b01010000; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01010110; c = 8'b01011101; // Expected: {'sum': 222, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01010110; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10110101; c = 8'b10011111; // Expected: {'sum': 71, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10110101; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00000101; c = 8'b10000111; // Expected: {'sum': 177, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00000101; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11100101; c = 8'b01111011; // Expected: {'sum': 104, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11100101; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10011000; c = 8'b10010100; // Expected: {'sum': 123, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10011000; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b00001010; c = 8'b11100010; // Expected: {'sum': 111, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b00001010; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01111110; c = 8'b10111010; // Expected: {'sum': 24, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01111110; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11100111; c = 8'b11111011; // Expected: {'sum': 168, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11100111; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10001011; c = 8'b11000001; // Expected: {'sum': 164, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10001011; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b01110101; c = 8'b11000111; // Expected: {'sum': 31, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b01110101; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11011111; c = 8'b00010001; // Expected: {'sum': 74, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11011111; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00000010; c = 8'b11011100; // Expected: {'sum': 104, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00000010; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b01011101; c = 8'b10001000; // Expected: {'sum': 65, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b01011101; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10011111; c = 8'b10101010; // Expected: {'sum': 218, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10011111; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10110111; c = 8'b00100000; // Expected: {'sum': 249, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10110111; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01010111; c = 8'b01100001; // Expected: {'sum': 93, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01010111; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00101000; c = 8'b01001000; // Expected: {'sum': 36, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00101000; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b01010000; c = 8'b00000111; // Expected: {'sum': 42, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b01010000; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10100011; c = 8'b10100110; // Expected: {'sum': 165, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10100011; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b11010101; c = 8'b00000110; // Expected: {'sum': 244, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b11010101; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00110010; c = 8'b11110111; // Expected: {'sum': 214, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00110010; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00110000; c = 8'b10010001; // Expected: {'sum': 79, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00110000; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b00001010; c = 8'b10001001; // Expected: {'sum': 152, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b00001010; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b01001001; c = 8'b10010000; // Expected: {'sum': 195, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b01001001; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10111110; c = 8'b10111101; // Expected: {'sum': 101, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10111110; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11111000; c = 8'b11100000; // Expected: {'sum': 85, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11111000; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11011000; c = 8'b10011111; // Expected: {'sum': 54, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11011000; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10000001; c = 8'b01010010; // Expected: {'sum': 158, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10000001; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11110101; c = 8'b01111110; // Expected: {'sum': 201, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11110101; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b11011111; c = 8'b00010111; // Expected: {'sum': 33, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b11011111; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10110000; c = 8'b01010001; // Expected: {'sum': 8, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10110000; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10100001; c = 8'b11010011; // Expected: {'sum': 92, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10100001; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10010110; c = 8'b11001110; // Expected: {'sum': 96, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10010110; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00010010; c = 8'b01100101; // Expected: {'sum': 245, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00010010; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00011110; c = 8'b11011000; // Expected: {'sum': 118, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00011110; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10000110; c = 8'b00111010; // Expected: {'sum': 20, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10000110; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b01111110; c = 8'b11110010; // Expected: {'sum': 111, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b01111110; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11001101; c = 8'b11110010; // Expected: {'sum': 40, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11001101; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10001001; c = 8'b11010110; // Expected: {'sum': 99, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10001001; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01111011; c = 8'b11000101; // Expected: {'sum': 43, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01111011; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10001001; c = 8'b10101001; // Expected: {'sum': 71, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10001001; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11000000; c = 8'b00110110; // Expected: {'sum': 139, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11000000; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01100100; c = 8'b10111010; // Expected: {'sum': 209, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01100100; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00110001; c = 8'b11010010; // Expected: {'sum': 93, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00110001; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01111000; c = 8'b00110001; // Expected: {'sum': 85, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01111000; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11111001; c = 8'b10000111; // Expected: {'sum': 229, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11111001; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11011011; c = 8'b11111001; // Expected: {'sum': 45, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11011011; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11110111; c = 8'b10110101; // Expected: {'sum': 250, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11110111; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b10000011; c = 8'b00101110; // Expected: {'sum': 61, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b10000011; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01111100; c = 8'b00000100; // Expected: {'sum': 90, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01111100; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11001111; c = 8'b01110100; // Expected: {'sum': 1, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11001111; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10001110; c = 8'b01111111; // Expected: {'sum': 246, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10001110; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01100100; c = 8'b11001010; // Expected: {'sum': 158, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01100100; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b00000000; c = 8'b11100011; // Expected: {'sum': 62, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b00000000; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11101100; c = 8'b10101111; // Expected: {'sum': 15, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11101100; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b11001001; c = 8'b00000010; // Expected: {'sum': 230, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b11001001; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b11000000; c = 8'b10001011; // Expected: {'sum': 22, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b11000000; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00001001; c = 8'b01000001; // Expected: {'sum': 151, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00001001; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01100010; c = 8'b10100001; // Expected: {'sum': 88, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01100010; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11101110; c = 8'b10101000; // Expected: {'sum': 79, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11101110; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00101001; c = 8'b11010111; // Expected: {'sum': 178, 'carry': 77}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00101001; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00100111; c = 8'b11000101; // Expected: {'sum': 184, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00100111; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10101100; c = 8'b00011000; // Expected: {'sum': 31, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10101100; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11111011; c = 8'b10101101; // Expected: {'sum': 109, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11111011; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01110101; c = 8'b11010110; // Expected: {'sum': 231, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01110101; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10101110; c = 8'b01110001; // Expected: {'sum': 68, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10101110; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01011001; c = 8'b10010011; // Expected: {'sum': 39, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01011001; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00001011; c = 8'b10000101; // Expected: {'sum': 137, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00001011; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10100110; c = 8'b10111100; // Expected: {'sum': 68, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10100110; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b00000100; c = 8'b00011010; // Expected: {'sum': 185, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b00000100; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00100111; c = 8'b10010100; // Expected: {'sum': 179, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00100111; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10111010; c = 8'b01101111; // Expected: {'sum': 196, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10111010; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11111001; c = 8'b10100010; // Expected: {'sum': 142, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11111001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b00010101; c = 8'b00101000; // Expected: {'sum': 4, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b00010101; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11010010; c = 8'b00110101; // Expected: {'sum': 89, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11010010; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01000101; c = 8'b10000010; // Expected: {'sum': 53, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01000101; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b01010111; c = 8'b11000011; // Expected: {'sum': 161, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b01010111; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11000011; c = 8'b11010100; // Expected: {'sum': 201, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11000011; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b01001111; c = 8'b11111001; // Expected: {'sum': 119, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b01001111; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b00001011; c = 8'b10111100; // Expected: {'sum': 253, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b00001011; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10000001; c = 8'b01001100; // Expected: {'sum': 171, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10000001; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b10110110; c = 8'b11011110; // Expected: {'sum': 155, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b10110110; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b01100101; c = 8'b01101010; // Expected: {'sum': 245, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b01100101; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10101011; c = 8'b00000101; // Expected: {'sum': 60, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10101011; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b11011101; c = 8'b10111110; // Expected: {'sum': 129, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b11011101; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01001100; c = 8'b11000111; // Expected: {'sum': 91, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01001100; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01100001; c = 8'b00001011; // Expected: {'sum': 78, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01100001; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10000110; c = 8'b10110100; // Expected: {'sum': 55, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10000110; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10001010; c = 8'b11101000; // Expected: {'sum': 137, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10001010; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00011111; c = 8'b01011100; // Expected: {'sum': 189, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00011111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10100011; c = 8'b00001010; // Expected: {'sum': 124, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10100011; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01000111; c = 8'b00011000; // Expected: {'sum': 119, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01000111; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01111011; c = 8'b10010011; // Expected: {'sum': 126, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01111011; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00100101; c = 8'b11111101; // Expected: {'sum': 157, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00100101; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11111001; c = 8'b11111101; // Expected: {'sum': 8, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11111001; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10001100; c = 8'b10110111; // Expected: {'sum': 91, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10001100; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10010001; c = 8'b01010110; // Expected: {'sum': 226, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10010001; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01101000; c = 8'b11101001; // Expected: {'sum': 119, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01101000; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10001110; c = 8'b11100101; // Expected: {'sum': 228, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10001110; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01001111; c = 8'b01000001; // Expected: {'sum': 86, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01001111; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11100010; c = 8'b00000011; // Expected: {'sum': 108, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11100010; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b11010011; c = 8'b11001100; // Expected: {'sum': 73, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b11010011; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10011011; c = 8'b10010101; // Expected: {'sum': 108, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10011011; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10010001; c = 8'b01000000; // Expected: {'sum': 234, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10010001; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01101010; c = 8'b11101011; // Expected: {'sum': 203, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01101010; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10001001; c = 8'b00100010; // Expected: {'sum': 251, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10001001; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b00100110; c = 8'b10101011; // Expected: {'sum': 10, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b00100110; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00000010; c = 8'b10000101; // Expected: {'sum': 52, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00000010; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00101011; c = 8'b00100111; // Expected: {'sum': 230, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00101011; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b00010111; c = 8'b00001110; // Expected: {'sum': 210, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b00010111; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00100000; c = 8'b10101101; // Expected: {'sum': 207, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00100000; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01010110; c = 8'b01111110; // Expected: {'sum': 231, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01010110; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00000101; c = 8'b11111110; // Expected: {'sum': 232, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00000101; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11000100; c = 8'b11110010; // Expected: {'sum': 142, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11000100; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11001111; c = 8'b10101101; // Expected: {'sum': 143, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11001111; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00011100; c = 8'b00000101; // Expected: {'sum': 68, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00011100; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00111101; c = 8'b10101000; // Expected: {'sum': 12, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00111101; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b11111100; c = 8'b11101100; // Expected: {'sum': 2, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b11111100; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00110111; c = 8'b01100010; // Expected: {'sum': 168, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00110111; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b11110101; c = 8'b01111010; // Expected: {'sum': 84, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b11110101; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10111111; c = 8'b00000111; // Expected: {'sum': 194, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10111111; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01010111; c = 8'b11110111; // Expected: {'sum': 83, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01010111; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10101010; c = 8'b01001100; // Expected: {'sum': 82, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10101010; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11101101; c = 8'b11100010; // Expected: {'sum': 86, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11101101; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10111110; c = 8'b00011000; // Expected: {'sum': 190, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10111110; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01011011; c = 8'b01111010; // Expected: {'sum': 17, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01011011; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11110011; c = 8'b00110111; // Expected: {'sum': 124, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11110011; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11100111; c = 8'b00111000; // Expected: {'sum': 70, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11100111; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b00101000; c = 8'b10011110; // Expected: {'sum': 228, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b00101000; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11011010; c = 8'b10010101; // Expected: {'sum': 164, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11011010; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10110100; c = 8'b10001110; // Expected: {'sum': 219, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10110100; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11000110; c = 8'b11110011; // Expected: {'sum': 114, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11000110; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10101101; c = 8'b11011000; // Expected: {'sum': 169, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10101101; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11001011; c = 8'b01011110; // Expected: {'sum': 61, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11001011; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10010101; c = 8'b10001001; // Expected: {'sum': 5, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10010101; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01000111; c = 8'b10010100; // Expected: {'sum': 144, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01000111; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00010010; c = 8'b00111010; // Expected: {'sum': 5, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00010010; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11101010; c = 8'b11010011; // Expected: {'sum': 220, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11101010; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10110110; c = 8'b10110001; // Expected: {'sum': 179, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10110110; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b00010000; c = 8'b01111100; // Expected: {'sum': 194, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b00010000; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b01001110; c = 8'b00110101; // Expected: {'sum': 165, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b01001110; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11011101; c = 8'b00011011; // Expected: {'sum': 114, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11011101; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01010100; c = 8'b00001010; // Expected: {'sum': 194, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01010100; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b00101111; c = 8'b00110010; // Expected: {'sum': 15, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b00101111; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b01010100; c = 8'b01001101; // Expected: {'sum': 147, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b01010100; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b11010000; c = 8'b11000000; // Expected: {'sum': 178, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b11010000; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b10101010; c = 8'b10010010; // Expected: {'sum': 131, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b10101010; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10010110; c = 8'b10010111; // Expected: {'sum': 224, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10010110; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b00100001; c = 8'b11000000; // Expected: {'sum': 94, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b00100001; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b00010011; c = 8'b01001010; // Expected: {'sum': 13, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b00010011; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00111101; c = 8'b01111111; // Expected: {'sum': 14, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00111101; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00001111; c = 8'b10000101; // Expected: {'sum': 139, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00001111; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10110010; c = 8'b00100111; // Expected: {'sum': 109, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10110010; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11010011; c = 8'b10001010; // Expected: {'sum': 107, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11010011; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10000101; c = 8'b00001100; // Expected: {'sum': 47, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10000101; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00001001; c = 8'b00101110; // Expected: {'sum': 169, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00001001; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00111010; c = 8'b11000000; // Expected: {'sum': 230, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00111010; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10101001; c = 8'b10011111; // Expected: {'sum': 153, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10101001; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11101011; c = 8'b11111100; // Expected: {'sum': 198, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11101011; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b10000101; c = 8'b10000001; // Expected: {'sum': 184, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b10000101; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b01100100; c = 8'b10100111; // Expected: {'sum': 33, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b01100100; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00001010; c = 8'b00110000; // Expected: {'sum': 63, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00001010; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01101010; c = 8'b00011100; // Expected: {'sum': 151, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01101010; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b00011110; c = 8'b11001010; // Expected: {'sum': 174, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b00011110; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11100000; c = 8'b10001010; // Expected: {'sum': 186, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11100000; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00001010; c = 8'b10001101; // Expected: {'sum': 62, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00001010; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b00011001; c = 8'b01110000; // Expected: {'sum': 213, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b00011001; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01111010; c = 8'b10011100; // Expected: {'sum': 19, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01111010; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10101110; c = 8'b01000011; // Expected: {'sum': 43, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10101110; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11000001; c = 8'b10100111; // Expected: {'sum': 134, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11000001; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b11001000; c = 8'b00101010; // Expected: {'sum': 85, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b11001000; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10011100; c = 8'b01111011; // Expected: {'sum': 217, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10011100; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00110001; c = 8'b00000101; // Expected: {'sum': 181, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00110001; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01101101; c = 8'b10011100; // Expected: {'sum': 199, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01101101; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00101110; c = 8'b00001010; // Expected: {'sum': 243, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00101110; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b01000000; c = 8'b11110000; // Expected: {'sum': 158, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b01000000; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01101011; c = 8'b11010010; // Expected: {'sum': 24, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01101011; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11001100; c = 8'b01100111; // Expected: {'sum': 90, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11001100; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10100001; c = 8'b11011001; // Expected: {'sum': 137, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10100001; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11110010; c = 8'b11011111; // Expected: {'sum': 108, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11110010; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01011111; c = 8'b01100101; // Expected: {'sum': 102, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01011111; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11111011; c = 8'b00000101; // Expected: {'sum': 2, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11111011; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00110011; c = 8'b11000111; // Expected: {'sum': 25, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00110011; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11011111; c = 8'b11100111; // Expected: {'sum': 1, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11011111; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01011001; c = 8'b11010010; // Expected: {'sum': 86, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01011001; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10111011; c = 8'b01000111; // Expected: {'sum': 53, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10111011; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b10011110; c = 8'b01010111; // Expected: {'sum': 202, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b10011110; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01000000; c = 8'b01001000; // Expected: {'sum': 15, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01000000; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b10101110; c = 8'b00010000; // Expected: {'sum': 179, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b10101110; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11010001; c = 8'b11101011; // Expected: {'sum': 248, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11010001; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01000000; c = 8'b11010101; // Expected: {'sum': 167, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01000000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11011000; c = 8'b00000000; // Expected: {'sum': 148, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11011000; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b11000101; c = 8'b10101110; // Expected: {'sum': 132, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b11000101; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10110100; c = 8'b00111001; // Expected: {'sum': 48, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10110100; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10010111; c = 8'b10001001; // Expected: {'sum': 173, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10010111; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01010100; c = 8'b11011110; // Expected: {'sum': 107, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01010100; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00100011; c = 8'b10100111; // Expected: {'sum': 5, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00100011; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00000101; c = 8'b01001001; // Expected: {'sum': 37, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00000101; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11010101; c = 8'b01110001; // Expected: {'sum': 34, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11010101; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b01000110; c = 8'b01110111; // Expected: {'sum': 81, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b01000110; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00000100; c = 8'b11101110; // Expected: {'sum': 118, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00000100; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b11010101; c = 8'b11101111; // Expected: {'sum': 140, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b11010101; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b00011111; c = 8'b10010011; // Expected: {'sum': 108, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b00011111; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00001000; c = 8'b10000111; // Expected: {'sum': 54, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00001000; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10110001; c = 8'b10101111; // Expected: {'sum': 164, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10110001; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11000111; c = 8'b10011000; // Expected: {'sum': 10, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11000111; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01011001; c = 8'b10001010; // Expected: {'sum': 40, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01011001; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00000100; c = 8'b11011011; // Expected: {'sum': 246, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00000100; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00011111; c = 8'b00111010; // Expected: {'sum': 171, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00011111; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00100101; c = 8'b10100011; // Expected: {'sum': 194, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00100101; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10111010; c = 8'b10010101; // Expected: {'sum': 114, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10111010; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01000001; c = 8'b01111100; // Expected: {'sum': 185, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01000001; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01100111; c = 8'b10110010; // Expected: {'sum': 105, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01100111; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01000100; c = 8'b10010110; // Expected: {'sum': 54, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01000100; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00101110; c = 8'b11100111; // Expected: {'sum': 13, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00101110; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10010110; c = 8'b00111100; // Expected: {'sum': 2, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10010110; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01111111; c = 8'b11110000; // Expected: {'sum': 223, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01111111; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00011110; c = 8'b01111011; // Expected: {'sum': 16, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00011110; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b01000010; c = 8'b10000010; // Expected: {'sum': 96, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b01000010; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b00110110; c = 8'b00011001; // Expected: {'sum': 136, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b00110110; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11111110; c = 8'b10000000; // Expected: {'sum': 88, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11111110; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11111110; c = 8'b01111010; // Expected: {'sum': 2, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11111110; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11110011; c = 8'b10011000; // Expected: {'sum': 115, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11110011; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10111000; c = 8'b01111000; // Expected: {'sum': 32, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10111000; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10111010; c = 8'b01111001; // Expected: {'sum': 19, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10111010; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b11100010; c = 8'b10001111; // Expected: {'sum': 130, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b11100010; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01001011; c = 8'b10010000; // Expected: {'sum': 200, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01001011; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10111001; c = 8'b11010111; // Expected: {'sum': 208, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10111001; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11011110; c = 8'b11101011; // Expected: {'sum': 61, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11011110; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01111000; c = 8'b01110010; // Expected: {'sum': 138, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01111000; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10101111; c = 8'b10010111; // Expected: {'sum': 240, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10101111; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b11010010; c = 8'b01000111; // Expected: {'sum': 34, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b11010010; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b01000001; c = 8'b11111000; // Expected: {'sum': 187, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b01000001; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01110000; c = 8'b01000011; // Expected: {'sum': 161, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01110000; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b01100101; c = 8'b01000101; // Expected: {'sum': 63, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b01100101; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b00011010; c = 8'b10011111; // Expected: {'sum': 134, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b00011010; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00010011; c = 8'b11000111; // Expected: {'sum': 68, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00010011; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01011111; c = 8'b01101100; // Expected: {'sum': 222, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01011111; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b01001001; c = 8'b10011011; // Expected: {'sum': 19, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b01001001; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b11101101; c = 8'b01000000; // Expected: {'sum': 15, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b11101101; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11111101; c = 8'b11010001; // Expected: {'sum': 173, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11111101; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11001100; c = 8'b10110001; // Expected: {'sum': 117, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11001100; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b01111011; c = 8'b10011011; // Expected: {'sum': 26, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b01111011; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b11000000; c = 8'b01001001; // Expected: {'sum': 137, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b11000000; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01101100; c = 8'b10111100; // Expected: {'sum': 11, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01101100; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10110101; c = 8'b11000011; // Expected: {'sum': 16, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10110101; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01101100; c = 8'b00011010; // Expected: {'sum': 193, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01101100; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00111011; c = 8'b01011000; // Expected: {'sum': 56, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00111011; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b11101101; c = 8'b11111000; // Expected: {'sum': 80, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b11101101; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00010011; c = 8'b00101110; // Expected: {'sum': 19, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00010011; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b00011111; c = 8'b11000011; // Expected: {'sum': 142, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b00011111; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11010011; c = 8'b01000001; // Expected: {'sum': 21, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11010011; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01010010; c = 8'b10100111; // Expected: {'sum': 46, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01010010; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10110010; c = 8'b01111011; // Expected: {'sum': 223, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10110010; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00011010; c = 8'b11010000; // Expected: {'sum': 134, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00011010; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b01100110; c = 8'b01000000; // Expected: {'sum': 29, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b01100110; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11000110; c = 8'b11111001; // Expected: {'sum': 89, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11000110; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10011001; c = 8'b01110111; // Expected: {'sum': 18, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10011001; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10011001; c = 8'b11100110; // Expected: {'sum': 216, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10011001; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b10101111; c = 8'b01001111; // Expected: {'sum': 238, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b10101111; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b00001111; c = 8'b00000010; // Expected: {'sum': 94, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b00001111; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b11111000; c = 8'b11100111; // Expected: {'sum': 56, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b11111000; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b10101000; c = 8'b01100100; // Expected: {'sum': 189, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b10101000; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b11111000; c = 8'b00011000; // Expected: {'sum': 205, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b11111000; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00011111; c = 8'b10000011; // Expected: {'sum': 217, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00011111; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b11001111; c = 8'b00011111; // Expected: {'sum': 147, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b11001111; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10111011; c = 8'b11010100; // Expected: {'sum': 46, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10111011; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10110010; c = 8'b00100101; // Expected: {'sum': 69, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10110010; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11100110; c = 8'b10101000; // Expected: {'sum': 142, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11100110; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10001101; c = 8'b10001110; // Expected: {'sum': 170, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10001101; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b11000100; c = 8'b11011110; // Expected: {'sum': 10, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b11000100; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10011111; c = 8'b10011001; // Expected: {'sum': 135, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10011111; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01001100; c = 8'b10100111; // Expected: {'sum': 3, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01001100; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11111011; c = 8'b01000110; // Expected: {'sum': 181, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11111011; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10110010; c = 8'b00101100; // Expected: {'sum': 39, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10110010; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11010111; c = 8'b11100000; // Expected: {'sum': 218, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11010111; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b00100000; c = 8'b10110110; // Expected: {'sum': 163, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b00100000; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b00010010; c = 8'b11010011; // Expected: {'sum': 252, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b00010010; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00001011; c = 8'b10011010; // Expected: {'sum': 97, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00001011; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b00011100; c = 8'b01110110; // Expected: {'sum': 86, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b00011100; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b11111101; c = 8'b10001111; // Expected: {'sum': 223, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b11111101; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01011100; c = 8'b00010000; // Expected: {'sum': 157, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01011100; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10101100; c = 8'b01111101; // Expected: {'sum': 2, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10101100; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b01101000; c = 8'b01010000; // Expected: {'sum': 13, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b01101000; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00001011; c = 8'b11000100; // Expected: {'sum': 33, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00001011; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01011000; c = 8'b00011001; // Expected: {'sum': 101, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01011000; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b10011011; c = 8'b01010111; // Expected: {'sum': 253, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b10011011; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11100110; c = 8'b10001100; // Expected: {'sum': 222, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11100110; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00100110; c = 8'b10100101; // Expected: {'sum': 237, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00100110; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b10011111; c = 8'b11001011; // Expected: {'sum': 95, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b10011111; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10110010; c = 8'b11110110; // Expected: {'sum': 8, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10110010; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00101110; c = 8'b01100111; // Expected: {'sum': 216, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00101110; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b00111111; c = 8'b11000000; // Expected: {'sum': 212, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b00111111; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00101110; c = 8'b10101000; // Expected: {'sum': 245, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00101110; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00110101; c = 8'b11000100; // Expected: {'sum': 81, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00110101; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10000000; c = 8'b01101010; // Expected: {'sum': 67, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10000000; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b00010101; c = 8'b10001110; // Expected: {'sum': 49, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b00010101; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b10100101; c = 8'b10101110; // Expected: {'sum': 126, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b10100101; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b01001100; c = 8'b11010001; // Expected: {'sum': 79, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b01001100; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b10000111; c = 8'b00111111; // Expected: {'sum': 3, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b10000111; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b00110000; c = 8'b10011000; // Expected: {'sum': 179, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b00110000; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01011100; c = 8'b00010110; // Expected: {'sum': 143, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01011100; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01101000; c = 8'b01000000; // Expected: {'sum': 118, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01101000; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11001010; c = 8'b10011011; // Expected: {'sum': 53, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11001010; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10101001; c = 8'b10111100; // Expected: {'sum': 101, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10101001; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00000100; c = 8'b11111001; // Expected: {'sum': 189, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00000100; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00101010; c = 8'b11101010; // Expected: {'sum': 194, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00101010; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01000110; c = 8'b10001100; // Expected: {'sum': 69, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01000110; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11010100; c = 8'b00000110; // Expected: {'sum': 51, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11010100; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10011111; c = 8'b01001111; // Expected: {'sum': 44, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10011111; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b11011100; c = 8'b10010001; // Expected: {'sum': 7, 'carry': 216}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b11011100; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00010011; c = 8'b10010100; // Expected: {'sum': 22, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00010011; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10110111; c = 8'b11001100; // Expected: {'sum': 193, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10110111; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00010011; c = 8'b00011110; // Expected: {'sum': 112, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00010011; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10111010; c = 8'b10110010; // Expected: {'sum': 139, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10111010; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10011001; c = 8'b11011001; // Expected: {'sum': 148, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10011001; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b00100111; c = 8'b00010000; // Expected: {'sum': 107, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b00100111; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b11101001; c = 8'b11001100; // Expected: {'sum': 227, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b11101001; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01011100; c = 8'b01100011; // Expected: {'sum': 131, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01011100; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11100100; c = 8'b10011100; // Expected: {'sum': 225, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11100100; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11101011; c = 8'b00110111; // Expected: {'sum': 60, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11101011; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01001101; c = 8'b01111111; // Expected: {'sum': 215, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01001101; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00110010; c = 8'b01001000; // Expected: {'sum': 105, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00110010; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b10000001; c = 8'b01011110; // Expected: {'sum': 33, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b10000001; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b11000011; c = 8'b00000000; // Expected: {'sum': 0, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b11000011; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11101101; c = 8'b11110101; // Expected: {'sum': 169, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11101101; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01100010; c = 8'b11100000; // Expected: {'sum': 184, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01100010; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10110101; c = 8'b10011010; // Expected: {'sum': 0, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10110101; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b10001000; c = 8'b00010001; // Expected: {'sum': 41, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b10001000; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b00101001; c = 8'b01110110; // Expected: {'sum': 71, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b00101001; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00000111; c = 8'b10110111; // Expected: {'sum': 216, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00000111; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11011100; c = 8'b01000111; // Expected: {'sum': 229, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11011100; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01011011; c = 8'b00000111; // Expected: {'sum': 229, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01011011; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01101111; c = 8'b10110111; // Expected: {'sum': 170, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01101111; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00001001; c = 8'b00010101; // Expected: {'sum': 167, 'carry': 25}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00001001; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11001100; c = 8'b10010001; // Expected: {'sum': 28, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11001100; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b11010011; c = 8'b01100001; // Expected: {'sum': 123, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b11010011; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00100100; c = 8'b01001101; // Expected: {'sum': 234, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00100100; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b11001000; c = 8'b11011001; // Expected: {'sum': 57, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b11001000; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b11000011; c = 8'b10111001; // Expected: {'sum': 93, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b11000011; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00110001; c = 8'b00011010; // Expected: {'sum': 142, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00110001; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10111011; c = 8'b01011111; // Expected: {'sum': 59, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10111011; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01000001; c = 8'b10011001; // Expected: {'sum': 166, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01000001; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10001100; c = 8'b01011011; // Expected: {'sum': 23, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10001100; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11001001; c = 8'b00000010; // Expected: {'sum': 216, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11001001; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00000111; c = 8'b00110011; // Expected: {'sum': 168, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00000111; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11111101; c = 8'b11111000; // Expected: {'sum': 149, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11111101; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01111011; c = 8'b11011101; // Expected: {'sum': 75, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01111011; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b11001110; c = 8'b10101111; // Expected: {'sum': 216, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b11001110; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01000011; c = 8'b11011100; // Expected: {'sum': 161, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01000011; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b11100111; c = 8'b10111100; // Expected: {'sum': 101, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b11100111; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01110000; c = 8'b00111011; // Expected: {'sum': 125, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01110000; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11111011; c = 8'b00101110; // Expected: {'sum': 13, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11111011; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10011110; c = 8'b00110111; // Expected: {'sum': 64, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10011110; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11010010; c = 8'b00011100; // Expected: {'sum': 133, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11010010; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11111010; c = 8'b10000101; // Expected: {'sum': 69, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11111010; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b11111111; c = 8'b01010011; // Expected: {'sum': 170, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b11111111; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00101110; c = 8'b01111100; // Expected: {'sum': 31, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00101110; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01011001; c = 8'b00001000; // Expected: {'sum': 238, 'carry': 25}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01011001; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b10111100; c = 8'b00000100; // Expected: {'sum': 51, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b10111100; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01111001; c = 8'b11110100; // Expected: {'sum': 138, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01111001; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b11111000; c = 8'b10101011; // Expected: {'sum': 149, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b11111000; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11010111; c = 8'b10010010; // Expected: {'sum': 237, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11010111; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b01011010; c = 8'b00011011; // Expected: {'sum': 243, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b01011010; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11111100; c = 8'b01111110; // Expected: {'sum': 129, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11111100; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b01011000; c = 8'b00111001; // Expected: {'sum': 32, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b01011000; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10011010; c = 8'b10110111; // Expected: {'sum': 162, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10011010; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01000010; c = 8'b00110001; // Expected: {'sum': 110, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01000010; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b00011101; c = 8'b10000101; // Expected: {'sum': 76, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b00011101; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01111010; c = 8'b00110111; // Expected: {'sum': 232, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01111010; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11100101; c = 8'b00100110; // Expected: {'sum': 136, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11100101; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11101011; c = 8'b11111011; // Expected: {'sum': 34, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11101011; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11110000; c = 8'b11111001; // Expected: {'sum': 123, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11110000; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01101001; c = 8'b11011010; // Expected: {'sum': 44, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01101001; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00000010; c = 8'b00110011; // Expected: {'sum': 64, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00000010; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00100100; c = 8'b01011000; // Expected: {'sum': 247, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00100100; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b11000110; c = 8'b11001001; // Expected: {'sum': 225, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b11000110; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10111001; c = 8'b00101000; // Expected: {'sum': 140, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10111001; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b10100000; c = 8'b01000001; // Expected: {'sum': 187, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b10100000; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b11000001; c = 8'b01000101; // Expected: {'sum': 77, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b11000001; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00001100; c = 8'b10101001; // Expected: {'sum': 21, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00001100; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01101011; c = 8'b00010010; // Expected: {'sum': 246, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01101011; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10011010; c = 8'b01010010; // Expected: {'sum': 113, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10011010; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00101010; c = 8'b11011010; // Expected: {'sum': 48, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00101010; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11000100; c = 8'b11110001; // Expected: {'sum': 123, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11000100; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10110111; c = 8'b10100000; // Expected: {'sum': 239, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10110111; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b11000001; c = 8'b11010001; // Expected: {'sum': 76, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b11000001; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00010000; c = 8'b01001110; // Expected: {'sum': 133, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00010000; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01100001; c = 8'b01000110; // Expected: {'sum': 199, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01100001; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00110010; c = 8'b00000101; // Expected: {'sum': 60, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00110010; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00010010; c = 8'b11001110; // Expected: {'sum': 255, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00010010; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10010111; c = 8'b00001010; // Expected: {'sum': 253, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10010111; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10111101; c = 8'b01111000; // Expected: {'sum': 199, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10111101; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11111101; c = 8'b01101001; // Expected: {'sum': 211, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11111101; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00111101; c = 8'b11000111; // Expected: {'sum': 15, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00111101; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b10000101; c = 8'b10101100; // Expected: {'sum': 202, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b10000101; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01001011; c = 8'b00110011; // Expected: {'sum': 200, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01001011; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b01010100; c = 8'b00011001; // Expected: {'sum': 84, 'carry': 25}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b01010100; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01111101; c = 8'b10001110; // Expected: {'sum': 175, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01111101; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00110000; c = 8'b00011111; // Expected: {'sum': 108, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00110000; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b10000100; c = 8'b11111000; // Expected: {'sum': 50, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b10000100; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11010001; c = 8'b10101101; // Expected: {'sum': 173, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11010001; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b01011111; c = 8'b11010111; // Expected: {'sum': 198, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b01011111; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00111111; c = 8'b11000010; // Expected: {'sum': 153, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00111111; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b01110011; c = 8'b10110001; // Expected: {'sum': 64, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b01110011; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10111011; c = 8'b00011011; // Expected: {'sum': 82, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10111011; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00000000; c = 8'b00000001; // Expected: {'sum': 169, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00000000; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b11001110; c = 8'b10000101; // Expected: {'sum': 185, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b11001110; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10001001; c = 8'b10010001; // Expected: {'sum': 26, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10001001; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11001001; c = 8'b01011100; // Expected: {'sum': 224, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11001001; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b11101000; c = 8'b00111000; // Expected: {'sum': 192, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b11101000; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10100111; c = 8'b10101011; // Expected: {'sum': 47, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10100111; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00010011; c = 8'b11001111; // Expected: {'sum': 219, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00010011; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11101010; c = 8'b11110111; // Expected: {'sum': 38, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11101010; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b00000000; c = 8'b01010001; // Expected: {'sum': 71, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b00000000; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00001001; c = 8'b11001110; // Expected: {'sum': 202, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00001001; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b10100001; c = 8'b00101000; // Expected: {'sum': 237, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b10100001; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01000101; c = 8'b00110100; // Expected: {'sum': 57, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01000101; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01110111; c = 8'b00001001; // Expected: {'sum': 233, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01110111; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01011100; c = 8'b10111111; // Expected: {'sum': 104, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01011100; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00110111; c = 8'b01101010; // Expected: {'sum': 159, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00110111; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b11101100; c = 8'b00001010; // Expected: {'sum': 14, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b11101100; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b01011000; c = 8'b11001100; // Expected: {'sum': 142, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b01011000; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11011000; c = 8'b01100011; // Expected: {'sum': 64, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11011000; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b01010111; c = 8'b01101111; // Expected: {'sum': 254, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b01010111; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11010011; c = 8'b00011111; // Expected: {'sum': 56, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11010011; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01111000; c = 8'b00011111; // Expected: {'sum': 208, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01111000; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10101011; c = 8'b01000010; // Expected: {'sum': 243, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10101011; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10010010; c = 8'b10001011; // Expected: {'sum': 33, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10010010; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00011100; c = 8'b01100010; // Expected: {'sum': 91, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00011100; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b11110010; c = 8'b01110100; // Expected: {'sum': 182, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b11110010; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00001110; c = 8'b01110011; // Expected: {'sum': 97, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00001110; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b00001111; c = 8'b10011110; // Expected: {'sum': 170, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b00001111; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00100011; c = 8'b10011001; // Expected: {'sum': 17, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00100011; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b00001101; c = 8'b01010101; // Expected: {'sum': 237, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b00001101; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11100111; c = 8'b10100101; // Expected: {'sum': 22, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11100111; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b11100011; c = 8'b00001101; // Expected: {'sum': 135, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b11100011; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10100010; c = 8'b10000110; // Expected: {'sum': 105, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10100010; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01100000; c = 8'b11011011; // Expected: {'sum': 35, 'carry': 216}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01100000; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00111000; c = 8'b10101010; // Expected: {'sum': 37, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00111000; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01011000; c = 8'b11010111; // Expected: {'sum': 187, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01011000; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00010001; c = 8'b00010111; // Expected: {'sum': 243, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00010001; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01000001; c = 8'b01010111; // Expected: {'sum': 167, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01000001; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00001111; c = 8'b11110010; // Expected: {'sum': 127, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00001111; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00000001; c = 8'b00011101; // Expected: {'sum': 40, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00000001; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00011011; c = 8'b10100110; // Expected: {'sum': 242, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00011011; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11000101; c = 8'b10001100; // Expected: {'sum': 142, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11000101; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00111101; c = 8'b01001100; // Expected: {'sum': 189, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00111101; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11111101; c = 8'b11101111; // Expected: {'sum': 69, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11111101; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b10011100; c = 8'b10011111; // Expected: {'sum': 36, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b10011100; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11010110; c = 8'b11000001; // Expected: {'sum': 46, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11010110; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10000011; c = 8'b00100001; // Expected: {'sum': 101, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10000011; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01101010; c = 8'b10100010; // Expected: {'sum': 214, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01101010; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b11100010; c = 8'b10111100; // Expected: {'sum': 49, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b11100010; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01101001; c = 8'b11110010; // Expected: {'sum': 16, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01101001; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11001000; c = 8'b11101111; // Expected: {'sum': 162, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11001000; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11000110; c = 8'b01110101; // Expected: {'sum': 102, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11000110; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10001000; c = 8'b11010101; // Expected: {'sum': 12, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10001000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11111011; c = 8'b11011101; // Expected: {'sum': 84, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11111011; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00111010; c = 8'b00111011; // Expected: {'sum': 76, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00111010; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10000110; c = 8'b10110010; // Expected: {'sum': 253, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10000110; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01010100; c = 8'b10000101; // Expected: {'sum': 116, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01010100; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b11001111; c = 8'b11001000; // Expected: {'sum': 136, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b11001111; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b01001000; c = 8'b00110101; // Expected: {'sum': 64, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b01001000; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b01100111; c = 8'b00010101; // Expected: {'sum': 119, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b01100111; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11111010; c = 8'b01010010; // Expected: {'sum': 18, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11111010; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11110010; c = 8'b00101000; // Expected: {'sum': 205, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11110010; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11111110; c = 8'b10111000; // Expected: {'sum': 1, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11111110; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10010010; c = 8'b10111000; // Expected: {'sum': 79, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10010010; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00000010; c = 8'b10101001; // Expected: {'sum': 174, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00000010; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10010000; c = 8'b00011100; // Expected: {'sum': 233, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10010000; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b01101110; c = 8'b11111011; // Expected: {'sum': 222, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b01101110; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00011111; c = 8'b10010101; // Expected: {'sum': 121, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00011111; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00001000; c = 8'b00010110; // Expected: {'sum': 170, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00001000; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b01001111; c = 8'b10100011; // Expected: {'sum': 36, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b01001111; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b10000110; c = 8'b00011010; // Expected: {'sum': 123, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b10000110; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10110010; c = 8'b10111011; // Expected: {'sum': 94, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10110010; c = 8'b10111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10000100; c = 8'b00111010; // Expected: {'sum': 220, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10000100; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b11010011; c = 8'b10011000; // Expected: {'sum': 168, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b11010011; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00000000; c = 8'b10111100; // Expected: {'sum': 180, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00000000; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b01000010; c = 8'b01100011; // Expected: {'sum': 92, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b01000010; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b11111101; c = 8'b00000101; // Expected: {'sum': 86, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b11111101; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b00000111; c = 8'b00010010; // Expected: {'sum': 73, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b00000111; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11010101; c = 8'b01100101; // Expected: {'sum': 156, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11010101; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11101000; c = 8'b01110110; // Expected: {'sum': 98, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11101000; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10010100; c = 8'b11111111; // Expected: {'sum': 77, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10010100; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b10010100; c = 8'b11001100; // Expected: {'sum': 30, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b10010100; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10000010; c = 8'b10010000; // Expected: {'sum': 166, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10000010; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10100110; c = 8'b11100001; // Expected: {'sum': 149, 'carry': 226}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10100110; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00001111; c = 8'b01101011; // Expected: {'sum': 39, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00001111; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01001000; c = 8'b11101011; // Expected: {'sum': 142, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01001000; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b11101011; c = 8'b11010100; // Expected: {'sum': 117, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b11101011; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b10000100; c = 8'b01100000; // Expected: {'sum': 37, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b10000100; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b11111100; c = 8'b01111100; // Expected: {'sum': 45, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b11111100; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b00101010; c = 8'b10000010; // Expected: {'sum': 224, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b00101010; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b01011111; c = 8'b10101000; // Expected: {'sum': 41, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b01011111; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10000100; c = 8'b10000100; // Expected: {'sum': 217, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10000100; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00111010; c = 8'b11101100; // Expected: {'sum': 128, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00111010; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b01100010; c = 8'b01110101; // Expected: {'sum': 161, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b01100010; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 663,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b11000001; c = 8'b01111101; // Expected: {'sum': 116, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b11000001; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 664,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b11001101; c = 8'b11000000; // Expected: {'sum': 227, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b11001101; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 665,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00100001; c = 8'b10110010; // Expected: {'sum': 212, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00100001; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 666,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11011110; c = 8'b00111001; // Expected: {'sum': 194, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11011110; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 667,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b11101011; c = 8'b11100011; // Expected: {'sum': 34, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b11101011; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 668,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10100101; c = 8'b01101100; // Expected: {'sum': 125, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10100101; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 669,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01111010; c = 8'b01101010; // Expected: {'sum': 175, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01111010; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 670,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00100011; c = 8'b11110111; // Expected: {'sum': 46, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00100011; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 671,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10010011; c = 8'b01001111; // Expected: {'sum': 135, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10010011; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 672,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01101000; c = 8'b00010010; // Expected: {'sum': 42, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01101000; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 673,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11110010; c = 8'b01111010; // Expected: {'sum': 252, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11110010; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 674,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00110110; c = 8'b11000001; // Expected: {'sum': 222, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00110110; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 675,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01000001; c = 8'b01100100; // Expected: {'sum': 121, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01000001; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 676,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00001001; c = 8'b00010111; // Expected: {'sum': 36, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00001001; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 677,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00011000; c = 8'b01111110; // Expected: {'sum': 120, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00011000; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 678,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10110100; c = 8'b11111001; // Expected: {'sum': 235, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10110100; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 679,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11101100; c = 8'b00101011; // Expected: {'sum': 221, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11101100; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 680,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10011010; c = 8'b10000000; // Expected: {'sum': 163, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10011010; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 681,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b10111111; c = 8'b01000101; // Expected: {'sum': 105, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b10111111; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 682,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b01011110; c = 8'b01111001; // Expected: {'sum': 135, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b01011110; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 683,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01101100; c = 8'b01111000; // Expected: {'sum': 136, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01101100; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 684,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10110000; c = 8'b01110011; // Expected: {'sum': 135, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10110000; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 685,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01001000; c = 8'b10101101; // Expected: {'sum': 57, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01001000; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 686,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01011110; c = 8'b10000000; // Expected: {'sum': 130, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01011110; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 687,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00001010; c = 8'b01000110; // Expected: {'sum': 45, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00001010; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 688,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b10001001; c = 8'b00101111; // Expected: {'sum': 48, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b10001001; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 689,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10111100; c = 8'b01000000; // Expected: {'sum': 236, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10111100; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 690,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00010001; c = 8'b10001110; // Expected: {'sum': 96, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00010001; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 691,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01110111; c = 8'b00100001; // Expected: {'sum': 202, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01110111; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 692,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00001100; c = 8'b10110101; // Expected: {'sum': 154, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00001100; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 693,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b11110110; c = 8'b10000110; // Expected: {'sum': 12, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b11110110; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 694,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b00101011; c = 8'b11110101; // Expected: {'sum': 68, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b00101011; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 695,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11011010; c = 8'b01001011; // Expected: {'sum': 50, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11011010; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 696,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11100010; c = 8'b01110001; // Expected: {'sum': 186, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11100010; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 697,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01001111; c = 8'b00001011; // Expected: {'sum': 37, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01001111; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 698,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11001000; c = 8'b11100001; // Expected: {'sum': 62, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11001000; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 699,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b10010100; c = 8'b00110101; // Expected: {'sum': 146, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b10010100; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 700,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10010100; c = 8'b01110000; // Expected: {'sum': 174, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10010100; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 701,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01111111; c = 8'b01111010; // Expected: {'sum': 109, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01111111; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 702,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b10010000; c = 8'b01010000; // Expected: {'sum': 190, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b10010000; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 703,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11000011; c = 8'b00110011; // Expected: {'sum': 214, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11000011; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 704,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00011111; c = 8'b01001011; // Expected: {'sum': 141, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00011111; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 705,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b11100100; c = 8'b11011001; // Expected: {'sum': 97, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b11100100; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 706,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11000111; c = 8'b01101110; // Expected: {'sum': 92, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11000111; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 707,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11000101; c = 8'b00100110; // Expected: {'sum': 174, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11000101; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 708,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01110100; c = 8'b01101011; // Expected: {'sum': 167, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01110100; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 709,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b10100100; c = 8'b10110100; // Expected: {'sum': 88, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b10100100; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 710,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01110001; c = 8'b00010100; // Expected: {'sum': 189, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01110001; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 711,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11001011; c = 8'b01100010; // Expected: {'sum': 221, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11001011; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 712,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01101101; c = 8'b01101001; // Expected: {'sum': 139, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01101101; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 713,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01010001; c = 8'b10010011; // Expected: {'sum': 25, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01010001; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 714,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b11010001; c = 8'b01001101; // Expected: {'sum': 86, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b11010001; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 715,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00010100; c = 8'b00111101; // Expected: {'sum': 35, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00010100; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 716,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b10011110; c = 8'b00000110; // Expected: {'sum': 143, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b10011110; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 717,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00010111; c = 8'b11110110; // Expected: {'sum': 135, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00010111; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 718,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b11010010; c = 8'b01111010; // Expected: {'sum': 216, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b11010010; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 719,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00111010; c = 8'b01000011; // Expected: {'sum': 196, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00111010; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 720,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b10001011; c = 8'b11101100; // Expected: {'sum': 176, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b10001011; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 721,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01111101; c = 8'b01100110; // Expected: {'sum': 54, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01111101; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 722,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10111100; c = 8'b01110110; // Expected: {'sum': 78, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10111100; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 723,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00000000; c = 8'b11111011; // Expected: {'sum': 147, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00000000; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 724,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01010010; c = 8'b10111111; // Expected: {'sum': 175, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01010010; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 725,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b11010010; c = 8'b01001101; // Expected: {'sum': 101, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b11010010; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 726,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00101110; c = 8'b11110100; // Expected: {'sum': 32, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00101110; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 727,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10111001; c = 8'b00111111; // Expected: {'sum': 95, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10111001; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 728,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b11101101; c = 8'b10100000; // Expected: {'sum': 189, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b11101101; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 729,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01100010; c = 8'b11001010; // Expected: {'sum': 211, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01100010; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 730,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10001110; c = 8'b11101010; // Expected: {'sum': 169, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10001110; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 731,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b11011110; c = 8'b01111010; // Expected: {'sum': 235, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b11011110; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 732,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01111000; c = 8'b11001010; // Expected: {'sum': 90, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01111000; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 733,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11000000; c = 8'b00011010; // Expected: {'sum': 115, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11000000; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 734,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00110000; c = 8'b11011100; // Expected: {'sum': 13, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00110000; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 735,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b01011011; c = 8'b10111110; // Expected: {'sum': 243, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b01011011; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 736,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b11001001; c = 8'b10001111; // Expected: {'sum': 15, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b11001001; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 737,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01100000; c = 8'b00000111; // Expected: {'sum': 27, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01100000; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 738,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b11001011; c = 8'b10110010; // Expected: {'sum': 33, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b11001011; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 739,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10010011; c = 8'b11010011; // Expected: {'sum': 160, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10010011; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 740,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b00001001; c = 8'b01011011; // Expected: {'sum': 137, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b00001001; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 741,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b11101100; c = 8'b11100110; // Expected: {'sum': 52, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b11101100; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 742,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b00101000; c = 8'b11000100; // Expected: {'sum': 150, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b00101000; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 743,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11100001; c = 8'b11111101; // Expected: {'sum': 104, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11100001; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 744,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b01011010; c = 8'b11001100; // Expected: {'sum': 161, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b01011010; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 745,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11111110; c = 8'b01110100; // Expected: {'sum': 219, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11111110; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 746,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10010001; c = 8'b01000000; // Expected: {'sum': 84, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10010001; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 747,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b01110010; c = 8'b10000100; // Expected: {'sum': 182, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b01110010; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 748,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00001101; c = 8'b00100111; // Expected: {'sum': 217, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00001101; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 749,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00001000; c = 8'b11101000; // Expected: {'sum': 63, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00001000; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 750,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b10101101; c = 8'b11000101; // Expected: {'sum': 23, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b10101101; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 751,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b11111101; c = 8'b10110010; // Expected: {'sum': 234, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b11111101; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 752,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01110100; c = 8'b01111001; // Expected: {'sum': 132, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01110100; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 753,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10011000; c = 8'b00001101; // Expected: {'sum': 169, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10011000; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 754,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00000100; c = 8'b01101011; // Expected: {'sum': 136, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00000100; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 755,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01011110; c = 8'b10101101; // Expected: {'sum': 187, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01011110; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 756,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b00011111; c = 8'b00110001; // Expected: {'sum': 183, 'carry': 25}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b00011111; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 757,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b00111011; c = 8'b01111110; // Expected: {'sum': 75, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b00111011; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 758,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11111111; c = 8'b11011100; // Expected: {'sum': 98, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11111111; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 759,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01000110; c = 8'b01001010; // Expected: {'sum': 63, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01000110; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 760,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b10010010; c = 8'b11110001; // Expected: {'sum': 42, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b10010010; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 761,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10000110; c = 8'b10101101; // Expected: {'sum': 135, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10000110; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 762,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b11010101; c = 8'b01110011; // Expected: {'sum': 45, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b11010101; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 763,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00111001; c = 8'b00000001; // Expected: {'sum': 169, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00111001; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 764,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b11110010; c = 8'b00011110; // Expected: {'sum': 141, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b11110010; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 765,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10101110; c = 8'b10110111; // Expected: {'sum': 35, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10101110; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 766,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10001100; c = 8'b10010000; // Expected: {'sum': 162, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10001100; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 767,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b00000001; c = 8'b01000010; // Expected: {'sum': 142, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b00000001; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 768,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00001000; c = 8'b00101010; // Expected: {'sum': 93, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00001000; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 769,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11001000; c = 8'b00111001; // Expected: {'sum': 63, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11001000; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 770,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11010011; c = 8'b11000001; // Expected: {'sum': 202, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11010011; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 771,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01001101; c = 8'b10010100; // Expected: {'sum': 184, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01001101; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 772,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00011111; c = 8'b01100011; // Expected: {'sum': 150, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00011111; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 773,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b11100111; c = 8'b00100001; // Expected: {'sum': 175, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b11100111; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 774,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00010000; c = 8'b10001010; // Expected: {'sum': 107, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00010000; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 775,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00001010; c = 8'b11011111; // Expected: {'sum': 100, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00001010; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 776,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11101111; c = 8'b11011100; // Expected: {'sum': 144, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11101111; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 777,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01111100; c = 8'b01101110; // Expected: {'sum': 137, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01111100; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 778,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11111001; c = 8'b11110101; // Expected: {'sum': 200, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11111001; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 779,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b00001110; c = 8'b00000001; // Expected: {'sum': 200, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b00001110; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 780,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10111011; c = 8'b10010000; // Expected: {'sum': 115, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10111011; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 781,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01101111; c = 8'b10101011; // Expected: {'sum': 175, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01101111; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 782,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b00011001; c = 8'b10111000; // Expected: {'sum': 162, 'carry': 25}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b00011001; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 783,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10100101; c = 8'b10111100; // Expected: {'sum': 154, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10100101; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 784,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b00100111; c = 8'b00101010; // Expected: {'sum': 121, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b00100111; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 785,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b00010100; c = 8'b10100101; // Expected: {'sum': 150, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b00010100; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 786,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b00100010; c = 8'b10001101; // Expected: {'sum': 189, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b00100010; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 787,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b10011100; c = 8'b11010100; // Expected: {'sum': 95, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b10011100; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 788,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b00110101; c = 8'b00101110; // Expected: {'sum': 142, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b00110101; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 789,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01101011; c = 8'b11111111; // Expected: {'sum': 66, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01101011; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 790,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10110101; c = 8'b00100101; // Expected: {'sum': 51, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10110101; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 791,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00010001; c = 8'b01111011; // Expected: {'sum': 90, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00010001; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 792,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b01111011; c = 8'b10000111; // Expected: {'sum': 33, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b01111011; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 793,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00011011; c = 8'b01000011; // Expected: {'sum': 126, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00011011; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 794,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b10111100; c = 8'b10101110; // Expected: {'sum': 31, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b10111100; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 795,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01001100; c = 8'b11100001; // Expected: {'sum': 173, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01001100; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 796,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b01000101; c = 8'b01011110; // Expected: {'sum': 197, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b01000101; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 797,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b11100110; c = 8'b01100001; // Expected: {'sum': 73, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b11100110; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 798,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b01101100; c = 8'b10011001; // Expected: {'sum': 57, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b01101100; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 799,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b01011101; c = 8'b11111000; // Expected: {'sum': 209, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b01011101; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 800,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b11110100; c = 8'b11100011; // Expected: {'sum': 156, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b11110100; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 801,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b10100001; c = 8'b11101101; // Expected: {'sum': 62, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b10100001; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 802,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01001000; c = 8'b11110001; // Expected: {'sum': 225, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01001000; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 803,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10101011; c = 8'b10001101; // Expected: {'sum': 113, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10101011; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 804,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01110101; c = 8'b01010001; // Expected: {'sum': 64, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01110101; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 805,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00001011; c = 8'b11001011; // Expected: {'sum': 92, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00001011; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 806,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00110010; c = 8'b00010110; // Expected: {'sum': 153, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00110010; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 807,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b11101010; c = 8'b11001011; // Expected: {'sum': 170, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b11101010; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 808,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11000110; c = 8'b01010110; // Expected: {'sum': 143, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11000110; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 809,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b01101100; c = 8'b10010000; // Expected: {'sum': 92, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b01101100; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 810,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00110101; c = 8'b11011011; // Expected: {'sum': 17, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00110101; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 811,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00010110; c = 8'b11100010; // Expected: {'sum': 199, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00010110; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 812,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b11110110; c = 8'b11001111; // Expected: {'sum': 219, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b11110110; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 813,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00100011; c = 8'b00000011; // Expected: {'sum': 118, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00100011; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 814,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b01100110; c = 8'b11101010; // Expected: {'sum': 14, 'carry': 226}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b01100110; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 815,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01111110; c = 8'b10100000; // Expected: {'sum': 17, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01111110; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 816,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11010101; c = 8'b01000000; // Expected: {'sum': 177, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11010101; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 817,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01100101; c = 8'b00110101; // Expected: {'sum': 212, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01100101; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 818,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b01000111; c = 8'b00111101; // Expected: {'sum': 20, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b01000111; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 819,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01011111; c = 8'b01110011; // Expected: {'sum': 150, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01011111; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 820,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b10110011; c = 8'b11100001; // Expected: {'sum': 59, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b10110011; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 821,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b11111010; c = 8'b11001001; // Expected: {'sum': 133, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b11111010; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 822,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10111110; c = 8'b11000111; // Expected: {'sum': 75, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10111110; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 823,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01100001; c = 8'b01110110; // Expected: {'sum': 31, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01100001; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 824,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10000011; c = 8'b10010011; // Expected: {'sum': 235, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10000011; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 825,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b00101110; c = 8'b11101011; // Expected: {'sum': 139, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b00101110; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 826,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b10100111; c = 8'b10110001; // Expected: {'sum': 117, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b10100111; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 827,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10111010; c = 8'b10101101; // Expected: {'sum': 213, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10111010; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 828,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11111100; c = 8'b00111010; // Expected: {'sum': 165, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11111100; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 829,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10000111; c = 8'b11111010; // Expected: {'sum': 180, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10000111; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 830,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b00101010; c = 8'b00100001; // Expected: {'sum': 85, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b00101010; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 831,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b01010100; c = 8'b00010111; // Expected: {'sum': 35, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b01010100; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 832,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11001010; c = 8'b00010010; // Expected: {'sum': 152, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11001010; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 833,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10101001; c = 8'b10000100; // Expected: {'sum': 221, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10101001; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 834,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01011101; c = 8'b11110100; // Expected: {'sum': 210, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01011101; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 835,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11011010; c = 8'b10100000; // Expected: {'sum': 76, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11011010; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 836,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01010111; c = 8'b10010100; // Expected: {'sum': 200, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01010111; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 837,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10000000; c = 8'b10000001; // Expected: {'sum': 142, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10000000; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 838,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01011101; c = 8'b01100010; // Expected: {'sum': 206, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01011101; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 839,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01000000; c = 8'b11101001; // Expected: {'sum': 242, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01000000; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 840,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11011010; c = 8'b11001100; // Expected: {'sum': 50, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11011010; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 841,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b10000111; c = 8'b01001000; // Expected: {'sum': 144, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b10000111; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 842,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b10101111; c = 8'b01111110; // Expected: {'sum': 251, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b10101111; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 843,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10011010; c = 8'b10100111; // Expected: {'sum': 213, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10011010; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 844,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10010100; c = 8'b01010011; // Expected: {'sum': 150, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10010100; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 845,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10010100; c = 8'b00001110; // Expected: {'sum': 45, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10010100; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 846,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10010110; c = 8'b01101101; // Expected: {'sum': 63, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10010110; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 847,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00011110; c = 8'b01110000; // Expected: {'sum': 143, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00011110; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 848,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b01000111; c = 8'b10111100; // Expected: {'sum': 130, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b01000111; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 849,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10001011; c = 8'b11011001; // Expected: {'sum': 25, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10001011; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 850,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10110100; c = 8'b10100011; // Expected: {'sum': 15, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10110100; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 851,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11010110; c = 8'b11011001; // Expected: {'sum': 217, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11010110; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 852,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01011011; c = 8'b01110001; // Expected: {'sum': 165, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01011011; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 853,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b11010010; c = 8'b01011111; // Expected: {'sum': 44, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b11010010; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 854,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b11111100; c = 8'b11010111; // Expected: {'sum': 74, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b11111100; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 855,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01000001; c = 8'b00000001; // Expected: {'sum': 169, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01000001; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 856,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01001101; c = 8'b10110100; // Expected: {'sum': 116, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01001101; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 857,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10100111; c = 8'b01000110; // Expected: {'sum': 188, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10100111; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 858,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b11010111; c = 8'b10101110; // Expected: {'sum': 198, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b11010111; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 859,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10101010; c = 8'b11110011; // Expected: {'sum': 24, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10101010; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 860,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b01011010; c = 8'b11110010; // Expected: {'sum': 157, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b01011010; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 861,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10011110; c = 8'b01001100; // Expected: {'sum': 216, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10011110; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 862,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b00000100; c = 8'b00001000; // Expected: {'sum': 102, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b00000100; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 863,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10000101; c = 8'b00001001; // Expected: {'sum': 15, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10000101; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 864,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11100111; c = 8'b00011110; // Expected: {'sum': 130, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11100111; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 865,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b11001101; c = 8'b00011110; // Expected: {'sum': 76, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b11001101; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 866,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01111101; c = 8'b10001010; // Expected: {'sum': 213, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01111101; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 867,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01101110; c = 8'b11111100; // Expected: {'sum': 174, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01101110; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 868,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01001101; c = 8'b01000110; // Expected: {'sum': 79, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01001101; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 869,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01101110; c = 8'b10111000; // Expected: {'sum': 63, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01101110; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 870,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b11111000; c = 8'b11101110; // Expected: {'sum': 171, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b11111000; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 871,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b01101011; c = 8'b01111100; // Expected: {'sum': 144, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b01101011; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 872,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11000111; c = 8'b11010001; // Expected: {'sum': 231, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11000111; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 873,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00011001; c = 8'b00110000; // Expected: {'sum': 90, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00011001; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 874,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b01000100; c = 8'b11000110; // Expected: {'sum': 160, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b01000100; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 875,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00000101; c = 8'b11001110; // Expected: {'sum': 139, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00000101; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 876,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01111010; c = 8'b10101011; // Expected: {'sum': 194, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01111010; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 877,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b11011111; c = 8'b00111011; // Expected: {'sum': 100, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b11011111; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 878,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b01111011; c = 8'b11010100; // Expected: {'sum': 64, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b01111011; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 879,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01111100; c = 8'b01110010; // Expected: {'sum': 185, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01111100; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 880,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10101000; c = 8'b00010011; // Expected: {'sum': 86, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10101000; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 881,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b10001010; c = 8'b01100001; // Expected: {'sum': 230, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b10001010; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 882,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00001000; c = 8'b01110101; // Expected: {'sum': 19, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00001000; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 883,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11011000; c = 8'b00010010; // Expected: {'sum': 191, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11011000; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 884,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00111110; c = 8'b00001010; // Expected: {'sum': 29, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00111110; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 885,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b01100001; c = 8'b01001111; // Expected: {'sum': 11, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b01100001; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 886,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00111100; c = 8'b01110100; // Expected: {'sum': 180, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00111100; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 887,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10001011; c = 8'b01110001; // Expected: {'sum': 172, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10001011; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 888,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01000000; c = 8'b11110011; // Expected: {'sum': 249, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01000000; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 889,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10010111; c = 8'b00111011; // Expected: {'sum': 181, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10010111; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 890,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b11110110; c = 8'b01110011; // Expected: {'sum': 133, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b11110110; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 891,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b00010111; c = 8'b10101101; // Expected: {'sum': 89, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b00010111; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 892,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00100011; c = 8'b11101111; // Expected: {'sum': 201, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00100011; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 893,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01010011; c = 8'b10100110; // Expected: {'sum': 117, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01010011; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 894,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11000110; c = 8'b00001011; // Expected: {'sum': 19, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11000110; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 895,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01101000; c = 8'b01101010; // Expected: {'sum': 105, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01101000; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 896,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11001001; c = 8'b00011111; // Expected: {'sum': 173, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11001001; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 897,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01011000; c = 8'b01001011; // Expected: {'sum': 123, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01011000; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 898,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b10110011; c = 8'b00000110; // Expected: {'sum': 201, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b10110011; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 899,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00111101; c = 8'b10101001; // Expected: {'sum': 252, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00111101; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 900,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01001011; c = 8'b01001110; // Expected: {'sum': 141, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01001011; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 901,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b10101000; c = 8'b01011111; // Expected: {'sum': 9, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b10101000; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 902,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b11011010; c = 8'b01010110; // Expected: {'sum': 77, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b11011010; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 903,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00010000; c = 8'b10011100; // Expected: {'sum': 44, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00010000; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 904,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b01001101; c = 8'b01110001; // Expected: {'sum': 85, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b01001101; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 905,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01101011; c = 8'b11101000; // Expected: {'sum': 135, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01101011; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 906,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00101010; c = 8'b00010011; // Expected: {'sum': 152, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00101010; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 907,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00101111; c = 8'b11010101; // Expected: {'sum': 58, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00101111; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 908,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11000010; c = 8'b00010101; // Expected: {'sum': 244, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11000010; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 909,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b00100111; c = 8'b01010001; // Expected: {'sum': 147, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b00100111; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 910,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b10110110; c = 8'b00011011; // Expected: {'sum': 8, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b10110110; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 911,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10001000; c = 8'b10000011; // Expected: {'sum': 79, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10001000; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 912,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10101101; c = 8'b00110111; // Expected: {'sum': 94, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10101101; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 913,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01101101; c = 8'b11101010; // Expected: {'sum': 196, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01101101; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 914,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00011110; c = 8'b01110111; // Expected: {'sum': 219, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00011110; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 915,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00110111; c = 8'b00110000; // Expected: {'sum': 172, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00110111; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 916,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01010101; c = 8'b00000101; // Expected: {'sum': 184, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01010101; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 917,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b01111000; c = 8'b10111101; // Expected: {'sum': 204, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b01111000; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 918,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b00100011; c = 8'b01010111; // Expected: {'sum': 128, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b00100011; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 919,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01111001; c = 8'b01110011; // Expected: {'sum': 52, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01111001; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 920,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10001101; c = 8'b10010100; // Expected: {'sum': 78, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10001101; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 921,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01011011; c = 8'b10101110; // Expected: {'sum': 222, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01011011; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 922,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b11001001; c = 8'b01010100; // Expected: {'sum': 205, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b11001001; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 923,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01001001; c = 8'b00011111; // Expected: {'sum': 69, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01001001; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 924,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00011111; c = 8'b11110010; // Expected: {'sum': 192, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00011111; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 925,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b11000101; c = 8'b11111100; // Expected: {'sum': 203, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b11000101; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 926,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00011000; c = 8'b10001011; // Expected: {'sum': 160, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00011000; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 927,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11101001; c = 8'b01101011; // Expected: {'sum': 83, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11101001; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 928,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b10010010; c = 8'b11001001; // Expected: {'sum': 215, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b10010010; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 929,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11001011; c = 8'b11001010; // Expected: {'sum': 191, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11001011; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 930,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01010010; c = 8'b00010011; // Expected: {'sum': 224, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01010010; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 931,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00011000; c = 8'b11000110; // Expected: {'sum': 51, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00011000; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 932,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00100110; c = 8'b01000011; // Expected: {'sum': 181, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00100110; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 933,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b01011111; c = 8'b10001010; // Expected: {'sum': 17, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b01011111; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 934,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00100001; c = 8'b10011111; // Expected: {'sum': 95, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00100001; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 935,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b10001010; c = 8'b01101110; // Expected: {'sum': 48, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b10001010; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 936,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b01111100; c = 8'b11101010; // Expected: {'sum': 144, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b01111100; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 937,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00010100; c = 8'b11111111; // Expected: {'sum': 15, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00010100; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 938,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b00010100; c = 8'b01111100; // Expected: {'sum': 67, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b00010100; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 939,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10001000; c = 8'b11011100; // Expected: {'sum': 10, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10001000; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 940,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b00100100; c = 8'b01111011; // Expected: {'sum': 6, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b00100100; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 941,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b11110001; c = 8'b01100111; // Expected: {'sum': 20, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b11110001; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 942,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b10100100; c = 8'b11100010; // Expected: {'sum': 198, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b10100100; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 943,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b10111000; c = 8'b10001101; // Expected: {'sum': 74, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b10111000; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 944,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10001010; c = 8'b01010101; // Expected: {'sum': 201, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10001010; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 945,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11100100; c = 8'b00100100; // Expected: {'sum': 88, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11100100; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 946,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01110101; c = 8'b01100100; // Expected: {'sum': 77, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01110101; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 947,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00111000; c = 8'b10000101; // Expected: {'sum': 181, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00111000; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 948,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b11000000; c = 8'b01100101; // Expected: {'sum': 141, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b11000000; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 949,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00111101; c = 8'b00101110; // Expected: {'sum': 239, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00111101; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 950,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00110001; c = 8'b00100111; // Expected: {'sum': 235, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00110001; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 951,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10000001; c = 8'b10101111; // Expected: {'sum': 152, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10000001; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 952,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01111001; c = 8'b00010101; // Expected: {'sum': 16, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01111001; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 953,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11011001; c = 8'b11010010; // Expected: {'sum': 116, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11011001; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 954,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10011011; c = 8'b00101000; // Expected: {'sum': 13, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10011011; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 955,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b00000110; c = 8'b00001000; // Expected: {'sum': 44, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b00000110; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 956,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b11100100; c = 8'b10100100; // Expected: {'sum': 58, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b11100100; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 957,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b10000001; c = 8'b01110110; // Expected: {'sum': 142, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b10000001; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 958,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b10000100; c = 8'b00100100; // Expected: {'sum': 136, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b10000100; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 959,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11110111; c = 8'b00100001; // Expected: {'sum': 104, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11110111; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 960,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11010100; c = 8'b10010010; // Expected: {'sum': 122, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11010100; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 961,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10000001; c = 8'b01100110; // Expected: {'sum': 37, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10000001; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 962,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00100100; c = 8'b11111011; // Expected: {'sum': 218, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00100100; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 963,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11101000; c = 8'b01100110; // Expected: {'sum': 93, 'carry': 226}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11101000; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 964,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b10110111; c = 8'b01000100; // Expected: {'sum': 160, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b10110111; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 965,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01010010; c = 8'b00001100; // Expected: {'sum': 52, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01010010; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 966,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00001011; c = 8'b01010000; // Expected: {'sum': 105, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00001011; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 967,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10001010; c = 8'b01101111; // Expected: {'sum': 43, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10001010; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 968,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01100110; c = 8'b01000011; // Expected: {'sum': 143, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01100110; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 969,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10011111; c = 8'b10001110; // Expected: {'sum': 164, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10011111; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 970,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b00000001; c = 8'b11111000; // Expected: {'sum': 198, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b00000001; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 971,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00110010; c = 8'b10011010; // Expected: {'sum': 67, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00110010; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 972,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00100001; c = 8'b11100000; // Expected: {'sum': 129, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00100001; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 973,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b00101111; c = 8'b11110000; // Expected: {'sum': 74, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b00101111; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 974,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11000010; c = 8'b00100110; // Expected: {'sum': 78, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11000010; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 975,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10101011; c = 8'b10011110; // Expected: {'sum': 36, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10101011; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 976,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b01111001; c = 8'b00001000; // Expected: {'sum': 204, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b01111001; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 977,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b11011111; c = 8'b01010001; // Expected: {'sum': 220, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b11011111; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 978,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00011100; c = 8'b00101100; // Expected: {'sum': 61, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00011100; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 979,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00011100; c = 8'b01001111; // Expected: {'sum': 162, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00011100; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 980,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11111010; c = 8'b10110100; // Expected: {'sum': 42, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11111010; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 981,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11110100; c = 8'b01101000; // Expected: {'sum': 132, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11110100; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 982,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01000000; c = 8'b11100100; // Expected: {'sum': 20, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01000000; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 983,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10111010; c = 8'b01000111; // Expected: {'sum': 105, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10111010; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 984,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11100000; c = 8'b00110000; // Expected: {'sum': 1, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11100000; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 985,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11001010; c = 8'b01111100; // Expected: {'sum': 21, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11001010; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 986,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11011111; c = 8'b11100001; // Expected: {'sum': 140, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11011111; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 987,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01111111; c = 8'b10111000; // Expected: {'sum': 244, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01111111; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 988,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11010011; c = 8'b11011010; // Expected: {'sum': 151, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11010011; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 989,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01110011; c = 8'b01110001; // Expected: {'sum': 169, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01110011; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 990,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01110011; c = 8'b01010010; // Expected: {'sum': 75, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01110011; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 991,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b11011010; c = 8'b00110000; // Expected: {'sum': 80, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b11011010; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 992,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b11010110; c = 8'b01001101; // Expected: {'sum': 171, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b11010110; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 993,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b01001001; c = 8'b01100100; // Expected: {'sum': 14, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b01001001; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 994,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01100001; c = 8'b01111111; // Expected: {'sum': 91, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01100001; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 995,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00010100; c = 8'b00011101; // Expected: {'sum': 39, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00010100; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 996,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00110001; c = 8'b10011100; // Expected: {'sum': 210, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00110001; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 997,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b00101001; c = 8'b11011100; // Expected: {'sum': 221, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b00101001; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 998,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10111111; c = 8'b01001000; // Expected: {'sum': 218, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10111111; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 999,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b00111011; c = 8'b01110110; // Expected: {'sum': 67, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b00111011; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1000,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b00000111; c = 8'b11111010; // Expected: {'sum': 188, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b00000111; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1001,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b01011100; c = 8'b11101110; // Expected: {'sum': 153, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b01011100; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1002,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b01100001; c = 8'b10101101; // Expected: {'sum': 56, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b01100001; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1003,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10101110; c = 8'b01000011; // Expected: {'sum': 46, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10101110; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1004,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b11001110; c = 8'b11011101; // Expected: {'sum': 223, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b11001110; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1005,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b11101101; c = 8'b00110000; // Expected: {'sum': 181, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b11101101; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1006,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11101110; c = 8'b10011011; // Expected: {'sum': 196, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11101110; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1007,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b00110110; c = 8'b00000001; // Expected: {'sum': 69, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b00110110; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1008,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00101000; c = 8'b00001100; // Expected: {'sum': 104, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00101000; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1009,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11000101; c = 8'b10000011; // Expected: {'sum': 212, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11000101; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1010,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00111011; c = 8'b11110010; // Expected: {'sum': 229, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00111011; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1011,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01101110; c = 8'b10010001; // Expected: {'sum': 197, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01101110; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1012,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00111111; c = 8'b11110010; // Expected: {'sum': 137, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00111111; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1013,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00010101; c = 8'b01000110; // Expected: {'sum': 49, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00010101; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1014,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00110001; c = 8'b01010000; // Expected: {'sum': 241, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00110001; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1015,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b00011111; c = 8'b11000110; // Expected: {'sum': 108, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b00011111; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1016,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b01110100; c = 8'b11001010; // Expected: {'sum': 131, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b01110100; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1017,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10001011; c = 8'b00111000; // Expected: {'sum': 69, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10001011; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1018,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b01110011; c = 8'b01011110; // Expected: {'sum': 254, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b01110011; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1019,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b01011000; c = 8'b00011000; // Expected: {'sum': 185, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b01011000; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1020,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b01101010; c = 8'b01101001; // Expected: {'sum': 254, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b01101010; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1021,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01011110; c = 8'b11100010; // Expected: {'sum': 23, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01011110; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1022,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01100011; c = 8'b10010001; // Expected: {'sum': 42, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01100011; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1023,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00101001; c = 8'b00000110; // Expected: {'sum': 185, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00101001; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1024,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b00100100; c = 8'b00101101; // Expected: {'sum': 85, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b00100100; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1025,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110011; c = 8'b10100101; // Expected: {'sum': 180, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110011; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1026,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11100001; c = 8'b10010010; // Expected: {'sum': 193, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11100001; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1027,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00101110; c = 8'b01100000; // Expected: {'sum': 19, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00101110; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1028,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00010010; c = 8'b00100010; // Expected: {'sum': 227, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00010010; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1029,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b11100110; c = 8'b11000110; // Expected: {'sum': 160, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b11100110; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1030,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b00011100; c = 8'b10111111; // Expected: {'sum': 96, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b00011100; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1031,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10010011; c = 8'b11101001; // Expected: {'sum': 98, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10010011; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1032,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11111001; c = 8'b10101010; // Expected: {'sum': 173, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11111001; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1033,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01111100; c = 8'b00111101; // Expected: {'sum': 190, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01111100; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1034,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00110010; c = 8'b11010110; // Expected: {'sum': 247, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00110010; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1035,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10111000; c = 8'b01101100; // Expected: {'sum': 35, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10111000; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1036,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11011100; c = 8'b00101001; // Expected: {'sum': 149, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11011100; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1037,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b01011001; c = 8'b00011011; // Expected: {'sum': 56, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b01011001; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1038,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b01100000; c = 8'b00010101; // Expected: {'sum': 137, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b01100000; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1039,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00000000; c = 8'b10100001; // Expected: {'sum': 182, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00000000; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1040,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b00100110; c = 8'b00110001; // Expected: {'sum': 7, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b00100110; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1041,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b01100001; c = 8'b01100110; // Expected: {'sum': 75, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b01100001; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1042,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10100001; c = 8'b01111100; // Expected: {'sum': 37, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10100001; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1043,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11011111; c = 8'b10100000; // Expected: {'sum': 242, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11011111; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1044,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11111100; c = 8'b01010100; // Expected: {'sum': 28, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11111100; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1045,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10101110; c = 8'b01111010; // Expected: {'sum': 77, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10101110; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1046,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b00100000; c = 8'b01010000; // Expected: {'sum': 164, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b00100000; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1047,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b01011110; c = 8'b00001110; // Expected: {'sum': 89, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b01011110; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1048,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b11101100; c = 8'b11100100; // Expected: {'sum': 226, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b11101100; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1049,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01011001; c = 8'b10111000; // Expected: {'sum': 185, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01011001; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1050,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b00010110; c = 8'b11010101; // Expected: {'sum': 44, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b00010110; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1051,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01111111; c = 8'b10000001; // Expected: {'sum': 62, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01111111; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1052,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00011010; c = 8'b00001111; // Expected: {'sum': 239, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00011010; c = 8'b00001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1053,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10100001; c = 8'b10110101; // Expected: {'sum': 249, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10100001; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1054,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00001110; c = 8'b11110011; // Expected: {'sum': 57, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00001110; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1055,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b11011100; c = 8'b11111101; // Expected: {'sum': 252, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b11011100; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1056,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00111011; c = 8'b01101010; // Expected: {'sum': 130, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00111011; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1057,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b00111110; c = 8'b10001011; // Expected: {'sum': 22, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b00111110; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1058,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01010111; c = 8'b01000000; // Expected: {'sum': 159, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01010111; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1059,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10101100; c = 8'b11001001; // Expected: {'sum': 236, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10101100; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1060,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11110100; c = 8'b10011110; // Expected: {'sum': 123, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11110100; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1061,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b00111111; c = 8'b00000010; // Expected: {'sum': 67, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b00111111; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1062,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b11000100; c = 8'b11100000; // Expected: {'sum': 217, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b11000100; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1063,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b01111111; c = 8'b01101111; // Expected: {'sum': 87, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b01111111; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1064,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b00010000; c = 8'b00001011; // Expected: {'sum': 159, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b00010000; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1065,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11010011; c = 8'b01010001; // Expected: {'sum': 92, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11010011; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1066,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00000110; c = 8'b01011100; // Expected: {'sum': 241, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00000110; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1067,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00111111; c = 8'b10111010; // Expected: {'sum': 103, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00111111; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1068,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10111011; c = 8'b00001001; // Expected: {'sum': 114, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10111011; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1069,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11111010; c = 8'b01011111; // Expected: {'sum': 17, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11111010; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1070,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b01010011; c = 8'b10001000; // Expected: {'sum': 59, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b01010011; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1071,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10100110; c = 8'b11001100; // Expected: {'sum': 87, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10100110; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1072,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b01100101; c = 8'b01011011; // Expected: {'sum': 121, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b01100101; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1073,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11110101; c = 8'b11110010; // Expected: {'sum': 52, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11110101; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1074,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b00100010; c = 8'b11000011; // Expected: {'sum': 7, 'carry': 226}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b00100010; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1075,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00111100; c = 8'b00100111; // Expected: {'sum': 238, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00111100; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1076,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b00001101; c = 8'b01110011; // Expected: {'sum': 97, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b00001101; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1077,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11001010; c = 8'b00000000; // Expected: {'sum': 105, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11001010; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1078,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b00111010; c = 8'b11110000; // Expected: {'sum': 109, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b00111010; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1079,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b01011111; c = 8'b00010010; // Expected: {'sum': 122, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b01011111; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1080,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b11100101; c = 8'b11111111; // Expected: {'sum': 181, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b11100101; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1081,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01001001; c = 8'b00100001; // Expected: {'sum': 155, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01001001; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1082,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b10101001; c = 8'b10010010; // Expected: {'sum': 25, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b10101001; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1083,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01010001; c = 8'b00010100; // Expected: {'sum': 124, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01010001; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1084,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11010111; c = 8'b01010111; // Expected: {'sum': 138, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11010111; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1085,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11111000; c = 8'b11011010; // Expected: {'sum': 40, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11111000; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1086,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b01010100; c = 8'b01101110; // Expected: {'sum': 40, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b01010100; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1087,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11011100; c = 8'b11111100; // Expected: {'sum': 149, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11011100; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1088,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00111011; c = 8'b00110101; // Expected: {'sum': 98, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00111011; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1089,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b10101101; c = 8'b01000111; // Expected: {'sum': 112, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b10101101; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1090,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b00110100; c = 8'b00001111; // Expected: {'sum': 174, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b00110100; c = 8'b00001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1091,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11101101; c = 8'b10001110; // Expected: {'sum': 163, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11101101; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1092,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11001101; c = 8'b10011110; // Expected: {'sum': 167, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11001101; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1093,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10010010; c = 8'b11010101; // Expected: {'sum': 220, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10010010; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1094,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b01000101; c = 8'b11010001; // Expected: {'sum': 105, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b01000101; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1095,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b00100000; c = 8'b10110101; // Expected: {'sum': 173, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b00100000; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1096,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b11111100; c = 8'b10010010; // Expected: {'sum': 153, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b11111100; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1097,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10111001; c = 8'b11010000; // Expected: {'sum': 160, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10111001; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1098,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10011110; c = 8'b10010111; // Expected: {'sum': 254, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10011110; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1099,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10010000; c = 8'b01110000; // Expected: {'sum': 114, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10010000; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00101010; c = 8'b11101101; // Expected: {'sum': 205, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00101010; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b10010100; c = 8'b11011100; // Expected: {'sum': 17, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b10010100; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b11111011; c = 8'b10100100; // Expected: {'sum': 232, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b11111011; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00100110; c = 8'b01001111; // Expected: {'sum': 219, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00100110; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b00111101; c = 8'b10100111; // Expected: {'sum': 56, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b00111101; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b10000110; c = 8'b00010000; // Expected: {'sum': 88, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b10000110; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10010101; c = 8'b10010000; // Expected: {'sum': 99, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10010101; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00100101; c = 8'b00101101; // Expected: {'sum': 191, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00100101; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b11110011; c = 8'b01011111; // Expected: {'sum': 239, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b11110011; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b00100110; c = 8'b11001010; // Expected: {'sum': 250, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b00100110; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b10001111; c = 8'b01111001; // Expected: {'sum': 87, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b10001111; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11000101; c = 8'b10110110; // Expected: {'sum': 147, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11000101; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b11100001; c = 8'b00011001; // Expected: {'sum': 232, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b11100001; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b11110001; c = 8'b00010001; // Expected: {'sum': 93, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b11110001; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00000101; c = 8'b00111110; // Expected: {'sum': 9, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00000101; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10111101; c = 8'b11011000; // Expected: {'sum': 32, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10111101; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01010100; c = 8'b00010101; // Expected: {'sum': 226, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01010100; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00000011; c = 8'b11111101; // Expected: {'sum': 222, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00000011; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00010101; c = 8'b01100101; // Expected: {'sum': 108, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00010101; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10011011; c = 8'b11001010; // Expected: {'sum': 109, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10011011; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01001011; c = 8'b11110100; // Expected: {'sum': 190, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01001011; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01111000; c = 8'b01100110; // Expected: {'sum': 229, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01111000; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11000001; c = 8'b10110010; // Expected: {'sum': 42, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11000001; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01010111; c = 8'b10000111; // Expected: {'sum': 26, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01010111; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11011001; c = 8'b00011000; // Expected: {'sum': 105, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11011001; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b01111000; c = 8'b10011110; // Expected: {'sum': 171, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b01111000; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11111101; c = 8'b10101011; // Expected: {'sum': 56, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11111101; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b01010000; c = 8'b00001100; // Expected: {'sum': 105, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b01010000; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b11000010; c = 8'b10000111; // Expected: {'sum': 22, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b11000010; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01110101; c = 8'b00110010; // Expected: {'sum': 235, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01110101; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01001100; c = 8'b10011101; // Expected: {'sum': 46, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01001100; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00010101; c = 8'b10001001; // Expected: {'sum': 57, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00010101; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b00011000; c = 8'b11001101; // Expected: {'sum': 85, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b00011000; c = 8'b11001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00001011; c = 8'b10111010; // Expected: {'sum': 66, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00001011; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01100011; c = 8'b10100000; // Expected: {'sum': 134, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01100011; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b01010100; c = 8'b10011101; // Expected: {'sum': 137, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b01010100; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11100011; c = 8'b11010001; // Expected: {'sum': 61, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11100011; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01000010; c = 8'b00110101; // Expected: {'sum': 231, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01000010; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10010000; c = 8'b00000111; // Expected: {'sum': 77, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10010000; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b10100101; c = 8'b00101100; // Expected: {'sum': 244, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b10100101; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b11001001; c = 8'b10001001; // Expected: {'sum': 189, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b11001001; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b10000101; c = 8'b01000111; // Expected: {'sum': 130, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b10000101; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01100010; c = 8'b11101000; // Expected: {'sum': 157, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01100010; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01010000; c = 8'b11111010; // Expected: {'sum': 41, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01010000; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10010111; c = 8'b01010100; // Expected: {'sum': 53, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10010111; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11110110; c = 8'b11110001; // Expected: {'sum': 86, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11110110; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10111100; c = 8'b10100100; // Expected: {'sum': 18, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10111100; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00101010; c = 8'b10110001; // Expected: {'sum': 183, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00101010; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11000100; c = 8'b01011101; // Expected: {'sum': 17, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11000100; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01101011; c = 8'b10111101; // Expected: {'sum': 35, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01101011; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11111001; c = 8'b00110111; // Expected: {'sum': 56, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11111001; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11110110; c = 8'b11110110; // Expected: {'sum': 158, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11110110; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11101011; c = 8'b01110000; // Expected: {'sum': 99, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11101011; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10011001; c = 8'b10100001; // Expected: {'sum': 152, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10011001; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10101011; c = 8'b01111111; // Expected: {'sum': 11, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10101011; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11101000; c = 8'b11001001; // Expected: {'sum': 117, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11101000; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00110000; c = 8'b11001110; // Expected: {'sum': 74, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00110000; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10001111; c = 8'b10001001; // Expected: {'sum': 237, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10001111; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10010100; c = 8'b00010111; // Expected: {'sum': 1, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10010100; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11110111; c = 8'b01100100; // Expected: {'sum': 87, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11110111; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01010111; c = 8'b10011110; // Expected: {'sum': 57, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01010111; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11010101; c = 8'b10101001; // Expected: {'sum': 109, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11010101; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b00111011; c = 8'b00101000; // Expected: {'sum': 231, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b00111011; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10001110; c = 8'b10110101; // Expected: {'sum': 45, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10001110; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b01101011; c = 8'b10010100; // Expected: {'sum': 143, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b01101011; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11001001; c = 8'b10100101; // Expected: {'sum': 17, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11001001; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b00111000; c = 8'b10110000; // Expected: {'sum': 149, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b00111000; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b01011011; c = 8'b00111110; // Expected: {'sum': 105, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b01011011; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11010110; c = 8'b10010110; // Expected: {'sum': 81, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11010110; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01101010; c = 8'b10100001; // Expected: {'sum': 189, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01101010; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10110000; c = 8'b10011110; // Expected: {'sum': 176, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10110000; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b11110010; c = 8'b00001100; // Expected: {'sum': 103, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b11110010; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b00101000; c = 8'b11111010; // Expected: {'sum': 240, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b00101000; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10010100; c = 8'b00110000; // Expected: {'sum': 2, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10010100; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b00111111; c = 8'b10110011; // Expected: {'sum': 225, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b00111111; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b01000000; c = 8'b10101100; // Expected: {'sum': 250, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b01000000; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01101111; c = 8'b00100110; // Expected: {'sum': 125, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01101111; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b00000111; c = 8'b11110010; // Expected: {'sum': 91, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b00000111; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10011111; c = 8'b11101110; // Expected: {'sum': 88, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10011111; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b00100001; c = 8'b01101010; // Expected: {'sum': 53, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b00100001; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b01111110; c = 8'b10101100; // Expected: {'sum': 231, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b01111110; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b11110010; c = 8'b10111000; // Expected: {'sum': 155, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b11110010; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b10001100; c = 8'b01000111; // Expected: {'sum': 145, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b10001100; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b11110011; c = 8'b11111101; // Expected: {'sum': 8, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b11110011; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01000100; c = 8'b11011110; // Expected: {'sum': 38, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01000100; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10011011; c = 8'b01100111; // Expected: {'sum': 173, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10011011; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b01101111; c = 8'b10101010; // Expected: {'sum': 49, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b01101111; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00011111; c = 8'b00011001; // Expected: {'sum': 157, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00011111; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00100000; c = 8'b01111100; // Expected: {'sum': 171, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00100000; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11011000; c = 8'b00000011; // Expected: {'sum': 94, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11011000; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00110000; c = 8'b01111101; // Expected: {'sum': 77, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00110000; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01101010; c = 8'b10010001; // Expected: {'sum': 74, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01101010; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00111000; c = 8'b10001011; // Expected: {'sum': 57, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00111000; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11101101; c = 8'b10010100; // Expected: {'sum': 122, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11101101; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00110111; c = 8'b01101000; // Expected: {'sum': 193, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00110111; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b01100001; c = 8'b01101010; // Expected: {'sum': 246, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b01100001; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01000101; c = 8'b10111011; // Expected: {'sum': 233, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01000101; c = 8'b10111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b10000100; c = 8'b00000110; // Expected: {'sum': 237, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b10000100; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11001100; c = 8'b11100011; // Expected: {'sum': 38, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11001100; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11110110; c = 8'b00111111; // Expected: {'sum': 56, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11110110; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10010000; c = 8'b10010001; // Expected: {'sum': 60, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10010000; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11010100; c = 8'b00100011; // Expected: {'sum': 174, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11010100; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00011010; c = 8'b00010010; // Expected: {'sum': 187, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00011010; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b00011100; c = 8'b11000111; // Expected: {'sum': 34, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b00011100; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b01010010; c = 8'b11001101; // Expected: {'sum': 83, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b01010010; c = 8'b11001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b01011110; c = 8'b11110010; // Expected: {'sum': 111, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b01011110; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00010111; c = 8'b11101111; // Expected: {'sum': 239, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00010111; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01111001; c = 8'b11101010; // Expected: {'sum': 125, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01111001; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11110001; c = 8'b01000110; // Expected: {'sum': 232, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11110001; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b00110100; c = 8'b11010100; // Expected: {'sum': 155, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b00110100; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01010110; c = 8'b01101011; // Expected: {'sum': 220, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01010110; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b01111100; c = 8'b10000001; // Expected: {'sum': 157, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b01111100; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00101110; c = 8'b11000011; // Expected: {'sum': 239, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00101110; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01010101; c = 8'b00000001; // Expected: {'sum': 129, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01010101; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01100100; c = 8'b11111010; // Expected: {'sum': 230, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01100100; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01010111; c = 8'b01110011; // Expected: {'sum': 212, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01010111; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11100110; c = 8'b10101010; // Expected: {'sum': 38, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11100110; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b00111010; c = 8'b01100001; // Expected: {'sum': 43, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b00111010; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11110100; c = 8'b11010010; // Expected: {'sum': 2, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11110100; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b00100001; c = 8'b00011011; // Expected: {'sum': 191, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b00100001; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00001010; c = 8'b01001000; // Expected: {'sum': 193, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00001010; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00101011; c = 8'b00110000; // Expected: {'sum': 147, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00101011; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b00011010; c = 8'b01000011; // Expected: {'sum': 229, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b00011010; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b10100010; c = 8'b00110000; // Expected: {'sum': 205, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b10100010; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b01011100; c = 8'b01000100; // Expected: {'sum': 239, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b01011100; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00001111; c = 8'b01010110; // Expected: {'sum': 179, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00001111; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01010111; c = 8'b01000101; // Expected: {'sum': 59, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01010111; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01010110; c = 8'b00100110; // Expected: {'sum': 169, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01010110; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b01101101; c = 8'b01111001; // Expected: {'sum': 227, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b01101101; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10001011; c = 8'b10010101; // Expected: {'sum': 114, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10001011; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00010001; c = 8'b01101010; // Expected: {'sum': 144, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00010001; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11011111; c = 8'b00111000; // Expected: {'sum': 31, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11011111; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11011010; c = 8'b10110111; // Expected: {'sum': 44, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11011010; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11100101; c = 8'b11111111; // Expected: {'sum': 150, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11100101; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00110100; c = 8'b00110110; // Expected: {'sum': 119, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00110100; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10111001; c = 8'b11011111; // Expected: {'sum': 62, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10111001; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11000111; c = 8'b01000010; // Expected: {'sum': 37, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11000111; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b11101101; c = 8'b10101000; // Expected: {'sum': 206, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b11101101; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b10110011; c = 8'b01011101; // Expected: {'sum': 113, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b10110011; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10100101; c = 8'b10111110; // Expected: {'sum': 179, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10100101; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b11001110; c = 8'b01110111; // Expected: {'sum': 160, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b11001110; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01000000; c = 8'b11100000; // Expected: {'sum': 106, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01000000; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 106, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11101011; c = 8'b11110001; // Expected: {'sum': 100, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11101011; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10110110; c = 8'b10100000; // Expected: {'sum': 28, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10110110; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b10100100; c = 8'b10111111; // Expected: {'sum': 177, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b10100100; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10010110; c = 8'b01010111; // Expected: {'sum': 84, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10010110; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11101010; c = 8'b11011010; // Expected: {'sum': 12, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11101010; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10110101; c = 8'b10011110; // Expected: {'sum': 207, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10110101; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b01110010; c = 8'b10011111; // Expected: {'sum': 95, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b01110010; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00011100; c = 8'b11011101; // Expected: {'sum': 123, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00011100; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00010001; c = 8'b00111011; // Expected: {'sum': 42, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00010001; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00111100; c = 8'b11011000; // Expected: {'sum': 194, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00111100; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b10010011; c = 8'b00001010; // Expected: {'sum': 152, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b10010011; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10001111; c = 8'b10000101; // Expected: {'sum': 252, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10001111; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00000000; c = 8'b00101011; // Expected: {'sum': 156, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00000000; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01110100; c = 8'b00000001; // Expected: {'sum': 117, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01110100; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11110011; c = 8'b01000010; // Expected: {'sum': 54, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11110011; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b11111000; c = 8'b11101101; // Expected: {'sum': 221, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b11111000; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01101011; c = 8'b00010011; // Expected: {'sum': 212, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01101011; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b00110001; c = 8'b11110000; // Expected: {'sum': 23, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b00110001; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01010101; c = 8'b11010001; // Expected: {'sum': 43, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01010101; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01100111; c = 8'b10110001; // Expected: {'sum': 82, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01100111; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00100010; c = 8'b11011010; // Expected: {'sum': 209, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00100010; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b10001110; c = 8'b10000000; // Expected: {'sum': 21, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b10001110; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b01000100; c = 8'b11000101; // Expected: {'sum': 146, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b01000100; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11010010; c = 8'b10111100; // Expected: {'sum': 187, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11010010; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00010110; c = 8'b10111100; // Expected: {'sum': 174, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00010110; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b11110111; c = 8'b01011011; // Expected: {'sum': 69, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b11110111; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b00101100; c = 8'b10111000; // Expected: {'sum': 196, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b00101100; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b11101100; c = 8'b10001011; // Expected: {'sum': 20, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b11101100; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00111001; c = 8'b01101110; // Expected: {'sum': 234, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00111001; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b01101111; c = 8'b01111001; // Expected: {'sum': 160, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b01101111; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10100110; c = 8'b00101110; // Expected: {'sum': 64, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10100110; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11011011; c = 8'b11000011; // Expected: {'sum': 117, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11011011; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01010001; c = 8'b00111011; // Expected: {'sum': 100, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01010001; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b11100110; c = 8'b00010001; // Expected: {'sum': 241, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b11100110; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00101011; c = 8'b00010100; // Expected: {'sum': 159, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00101011; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00001001; c = 8'b10111110; // Expected: {'sum': 169, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00001001; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00001100; c = 8'b00000011; // Expected: {'sum': 228, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00001100; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00110011; c = 8'b01011101; // Expected: {'sum': 225, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00110011; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b01111011; c = 8'b10000110; // Expected: {'sum': 3, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b01111011; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10110001; c = 8'b10001111; // Expected: {'sum': 210, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10110001; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01010001; c = 8'b10111111; // Expected: {'sum': 146, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01010001; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11110011; c = 8'b01010100; // Expected: {'sum': 94, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11110011; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b01011011; c = 8'b00110101; // Expected: {'sum': 186, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b01011011; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b01010000; c = 8'b10110011; // Expected: {'sum': 251, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b01010000; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b11010000; c = 8'b00010111; // Expected: {'sum': 126, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b11010000; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01111100; c = 8'b11011001; // Expected: {'sum': 222, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01111100; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10001111; c = 8'b01010101; // Expected: {'sum': 247, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10001111; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b00101100; c = 8'b11100100; // Expected: {'sum': 211, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b00101100; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01110111; c = 8'b11001110; // Expected: {'sum': 204, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01110111; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01001110; c = 8'b00101101; // Expected: {'sum': 22, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01001110; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11001001; c = 8'b11010001; // Expected: {'sum': 49, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11001001; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00101100; c = 8'b11111001; // Expected: {'sum': 132, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00101100; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01010011; c = 8'b11100010; // Expected: {'sum': 208, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01010011; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11100101; c = 8'b11001010; // Expected: {'sum': 212, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11100101; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11110100; c = 8'b01010100; // Expected: {'sum': 182, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11110100; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b10100010; c = 8'b00010000; // Expected: {'sum': 134, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b10100010; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11110000; c = 8'b00111000; // Expected: {'sum': 134, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11110000; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01010000; c = 8'b01101001; // Expected: {'sum': 177, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01010000; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01110011; c = 8'b00110110; // Expected: {'sum': 196, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01110011; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b11001001; c = 8'b11101101; // Expected: {'sum': 57, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b11001001; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00101011; c = 8'b01110101; // Expected: {'sum': 179, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00101011; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10001001; c = 8'b10010010; // Expected: {'sum': 209, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10001001; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01110100; c = 8'b01101010; // Expected: {'sum': 245, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01110100; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00011111; c = 8'b11111101; // Expected: {'sum': 180, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00011111; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b11011110; c = 8'b00111010; // Expected: {'sum': 201, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b11011110; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b00010000; c = 8'b00001001; // Expected: {'sum': 107, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b00010000; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00000100; c = 8'b11101010; // Expected: {'sum': 100, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00000100; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b11010010; c = 8'b10001001; // Expected: {'sum': 24, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b11010010; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b00001010; c = 8'b11111000; // Expected: {'sum': 36, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b00001010; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00001001; c = 8'b11101101; // Expected: {'sum': 199, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00001001; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00010010; c = 8'b01001011; // Expected: {'sum': 214, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00010010; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b10100000; c = 8'b01110001; // Expected: {'sum': 136, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b10100000; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10111111; c = 8'b01111010; // Expected: {'sum': 143, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10111111; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b11111010; c = 8'b10110000; // Expected: {'sum': 230, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b11111010; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10000110; c = 8'b11101100; // Expected: {'sum': 223, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10000110; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b01101011; c = 8'b01001000; // Expected: {'sum': 167, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b01101011; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00000000; c = 8'b10101000; // Expected: {'sum': 207, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00000000; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10000000; c = 8'b10000011; // Expected: {'sum': 247, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10000000; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01101001; c = 8'b11101101; // Expected: {'sum': 7, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01101001; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11000101; c = 8'b11000110; // Expected: {'sum': 195, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11000101; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00011010; c = 8'b11011101; // Expected: {'sum': 30, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00011010; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10000010; c = 8'b00010011; // Expected: {'sum': 136, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10000010; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11011111; c = 8'b01101001; // Expected: {'sum': 35, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11011111; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10010000; c = 8'b00111010; // Expected: {'sum': 210, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10010000; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b11010111; c = 8'b00110000; // Expected: {'sum': 100, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b11010111; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01000111; c = 8'b10010001; // Expected: {'sum': 174, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01000111; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01010100; c = 8'b10101100; // Expected: {'sum': 173, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01010100; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11111111; c = 8'b01010000; // Expected: {'sum': 227, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11111111; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00011000; c = 8'b10100101; // Expected: {'sum': 236, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00011000; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00110011; c = 8'b11111011; // Expected: {'sum': 105, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00110011; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b11100011; c = 8'b01101011; // Expected: {'sum': 81, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b11100011; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b01101110; c = 8'b11000111; // Expected: {'sum': 196, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b01101110; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00011001; c = 8'b00101100; // Expected: {'sum': 48, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00011001; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11110101; c = 8'b10101100; // Expected: {'sum': 24, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11110101; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11110111; c = 8'b10000010; // Expected: {'sum': 128, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11110111; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b10111100; c = 8'b10110111; // Expected: {'sum': 246, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b10111100; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10000011; c = 8'b00011011; // Expected: {'sum': 82, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10000011; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b00110001; c = 8'b01000001; // Expected: {'sum': 87, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b00110001; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b11110101; c = 8'b11101001; // Expected: {'sum': 121, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b11110101; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b00100011; c = 8'b01010011; // Expected: {'sum': 71, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b00100011; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b00000011; c = 8'b10100001; // Expected: {'sum': 207, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b00000011; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00011011; c = 8'b10010110; // Expected: {'sum': 17, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00011011; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01000000; c = 8'b00010000; // Expected: {'sum': 204, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01000000; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b11101100; c = 8'b01011110; // Expected: {'sum': 65, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b11101100; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00011110; c = 8'b01111110; // Expected: {'sum': 121, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00011110; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01011100; c = 8'b10011001; // Expected: {'sum': 48, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01011100; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b00011011; c = 8'b00100100; // Expected: {'sum': 75, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b00011011; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b00100111; c = 8'b01001000; // Expected: {'sum': 49, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b00100111; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b01110111; c = 8'b10110100; // Expected: {'sum': 125, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b01110111; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b00000110; c = 8'b01000000; // Expected: {'sum': 48, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b00000110; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01110111; c = 8'b00101111; // Expected: {'sum': 13, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01110111; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11100101; c = 8'b01110101; // Expected: {'sum': 153, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11100101; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b00000001; c = 8'b11110101; // Expected: {'sum': 90, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b00000001; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01111000; c = 8'b11100011; // Expected: {'sum': 117, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01111000; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00001000; c = 8'b10011011; // Expected: {'sum': 18, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00001000; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11001010; c = 8'b10011001; // Expected: {'sum': 141, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11001010; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b00010010; c = 8'b00100110; // Expected: {'sum': 236, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b00010010; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b10001101; c = 8'b00000010; // Expected: {'sum': 8, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b10001101; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11011101; c = 8'b00000001; // Expected: {'sum': 186, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11011101; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00111011; c = 8'b11110001; // Expected: {'sum': 191, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00111011; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00001100; c = 8'b01101001; // Expected: {'sum': 178, 'carry': 77}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00001100; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b00011010; c = 8'b10100111; // Expected: {'sum': 127, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b00011010; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01101101; c = 8'b00010100; // Expected: {'sum': 144, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01101101; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b10101110; c = 8'b01000011; // Expected: {'sum': 72, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b10101110; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00110000; c = 8'b00100110; // Expected: {'sum': 10, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00110000; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00010101; c = 8'b01011100; // Expected: {'sum': 228, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00010101; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01110101; c = 8'b00100000; // Expected: {'sum': 15, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01110101; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b11010000; c = 8'b10000001; // Expected: {'sum': 240, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b11010000; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01101101; c = 8'b01011010; // Expected: {'sum': 56, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01101101; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10110111; c = 8'b11011110; // Expected: {'sum': 215, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10110111; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11011101; c = 8'b10011101; // Expected: {'sum': 36, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11011101; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11000110; c = 8'b01011101; // Expected: {'sum': 234, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11000110; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10111010; c = 8'b11010011; // Expected: {'sum': 153, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10111010; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01111100; c = 8'b10010001; // Expected: {'sum': 87, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01111100; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01111001; c = 8'b10100110; // Expected: {'sum': 173, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01111001; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10111111; c = 8'b00100100; // Expected: {'sum': 215, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10111111; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00011111; c = 8'b00111101; // Expected: {'sum': 253, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00011111; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b00011001; c = 8'b01101100; // Expected: {'sum': 234, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b00011001; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01010100; c = 8'b00011100; // Expected: {'sum': 231, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01010100; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b10111011; c = 8'b11111010; // Expected: {'sum': 120, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b10111011; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10000001; c = 8'b01011001; // Expected: {'sum': 151, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10000001; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00111001; c = 8'b01001100; // Expected: {'sum': 32, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00111001; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00111000; c = 8'b10001011; // Expected: {'sum': 178, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00111000; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b10000101; c = 8'b10011000; // Expected: {'sum': 36, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b10000101; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b01010111; c = 8'b10010110; // Expected: {'sum': 38, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b01010111; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11101011; c = 8'b10001011; // Expected: {'sum': 176, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11101011; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b10101010; c = 8'b10110111; // Expected: {'sum': 114, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b10101010; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00011010; c = 8'b11110111; // Expected: {'sum': 17, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00011010; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00101000; c = 8'b01010010; // Expected: {'sum': 22, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00101000; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b10010001; c = 8'b11101001; // Expected: {'sum': 202, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b10010001; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11101100; c = 8'b10111100; // Expected: {'sum': 23, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11101100; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10010101; c = 8'b01110011; // Expected: {'sum': 98, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10010101; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00111110; c = 8'b10011001; // Expected: {'sum': 55, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00111110; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b01011010; c = 8'b01101011; // Expected: {'sum': 76, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b01011010; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b11100010; c = 8'b11000011; // Expected: {'sum': 49, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b11100010; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11100111; c = 8'b00110110; // Expected: {'sum': 101, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11100111; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10000011; c = 8'b00111110; // Expected: {'sum': 10, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10000011; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11000110; c = 8'b01000110; // Expected: {'sum': 217, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11000110; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b00011001; c = 8'b10100000; // Expected: {'sum': 132, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b00011001; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00001000; c = 8'b00110011; // Expected: {'sum': 93, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00001000; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01100000; c = 8'b10111110; // Expected: {'sum': 168, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01100000; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00001110; c = 8'b10100100; // Expected: {'sum': 168, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00001110; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b00000000; c = 8'b10011010; // Expected: {'sum': 133, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b00000000; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00110101; c = 8'b10010011; // Expected: {'sum': 143, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00110101; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10000101; c = 8'b11111001; // Expected: {'sum': 4, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10000101; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b11110010; c = 8'b01100000; // Expected: {'sum': 252, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b11110010; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10010110; c = 8'b00011011; // Expected: {'sum': 168, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10010110; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10110110; c = 8'b11110001; // Expected: {'sum': 179, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10110110; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b00101011; c = 8'b10110110; // Expected: {'sum': 88, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b00101011; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b10111111; c = 8'b10111101; // Expected: {'sum': 247, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b10111111; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10001001; c = 8'b01010011; // Expected: {'sum': 182, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10001001; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10111001; c = 8'b10000011; // Expected: {'sum': 137, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10111001; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10111101; c = 8'b00111101; // Expected: {'sum': 111, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10111101; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11011010; c = 8'b00100001; // Expected: {'sum': 175, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11011010; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10110110; c = 8'b11011000; // Expected: {'sum': 25, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10110110; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b01001100; c = 8'b00101010; // Expected: {'sum': 188, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b01001100; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01001010; c = 8'b01010010; // Expected: {'sum': 68, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01001010; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10100010; c = 8'b00010001; // Expected: {'sum': 82, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10100010; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b00100100; c = 8'b11100001; // Expected: {'sum': 146, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b00100100; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b01101001; c = 8'b11000111; // Expected: {'sum': 82, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b01101001; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b11111100; c = 8'b01110001; // Expected: {'sum': 141, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b11111100; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b01101100; c = 8'b11001111; // Expected: {'sum': 187, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b01101100; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00011101; c = 8'b01000101; // Expected: {'sum': 13, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00011101; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10110001; c = 8'b00110000; // Expected: {'sum': 135, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10110001; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01101100; c = 8'b01101010; // Expected: {'sum': 245, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01101100; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b01110010; c = 8'b10101101; // Expected: {'sum': 57, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b01110010; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b10111000; c = 8'b01111100; // Expected: {'sum': 134, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b10111000; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00110101; c = 8'b00000010; // Expected: {'sum': 119, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00110101; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b11000010; c = 8'b10111100; // Expected: {'sum': 248, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b11000010; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00000000; c = 8'b10010010; // Expected: {'sum': 92, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00000000; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b00011000; c = 8'b10001000; // Expected: {'sum': 150, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b00011000; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b01110100; c = 8'b11001000; // Expected: {'sum': 54, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b01110100; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b01000100; c = 8'b00001100; // Expected: {'sum': 234, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b01000100; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11001110; c = 8'b01011001; // Expected: {'sum': 55, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11001110; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10100111; c = 8'b01011001; // Expected: {'sum': 94, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10100111; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b00010100; c = 8'b11110010; // Expected: {'sum': 168, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b00010100; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10101100; c = 8'b10001010; // Expected: {'sum': 64, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10101100; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b10100001; c = 8'b00101001; // Expected: {'sum': 164, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b10100001; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00100000; c = 8'b01000000; // Expected: {'sum': 214, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00100000; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b00011011; c = 8'b00001011; // Expected: {'sum': 153, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b00011011; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b11010110; c = 8'b10100000; // Expected: {'sum': 253, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b11010110; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11111110; c = 8'b01101100; // Expected: {'sum': 77, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11111110; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110001; c = 8'b11111000; // Expected: {'sum': 235, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110001; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11111000; c = 8'b00110100; // Expected: {'sum': 92, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11111000; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b00100010; c = 8'b01001110; // Expected: {'sum': 224, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b00100010; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01010000; c = 8'b10101000; // Expected: {'sum': 164, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01010000; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b10011010; c = 8'b11101011; // Expected: {'sum': 30, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b10011010; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11111001; c = 8'b01011111; // Expected: {'sum': 62, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11111001; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11110010; c = 8'b11110010; // Expected: {'sum': 254, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11110010; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10001110; c = 8'b01010110; // Expected: {'sum': 48, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10001110; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11001000; c = 8'b10111010; // Expected: {'sum': 20, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11001000; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00011011; c = 8'b00111000; // Expected: {'sum': 212, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00011011; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00000011; c = 8'b00101100; // Expected: {'sum': 160, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00000011; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11100100; c = 8'b10010101; // Expected: {'sum': 141, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11100100; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b00111001; c = 8'b10111100; // Expected: {'sum': 145, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b00111001; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00111101; c = 8'b10111010; // Expected: {'sum': 229, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00111101; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11010011; c = 8'b10010000; // Expected: {'sum': 80, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11010011; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b11111010; c = 8'b11010110; // Expected: {'sum': 128, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b11111010; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10000100; c = 8'b10000111; // Expected: {'sum': 171, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10000100; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10111100; c = 8'b00110100; // Expected: {'sum': 145, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10111100; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00111100; c = 8'b00001111; // Expected: {'sum': 68, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00111100; c = 8'b00001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b01101110; c = 8'b01100101; // Expected: {'sum': 69, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b01101110; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10001111; c = 8'b01100100; // Expected: {'sum': 76, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10001111; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b11100101; c = 8'b11000101; // Expected: {'sum': 97, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b11100101; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01110111; c = 8'b10011101; // Expected: {'sum': 228, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01110111; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b01011101; c = 8'b01101001; // Expected: {'sum': 174, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b01011101; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b10001101; c = 8'b01110000; // Expected: {'sum': 204, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b10001101; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10010110; c = 8'b11010001; // Expected: {'sum': 136, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10010110; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b01100001; c = 8'b00010001; // Expected: {'sum': 56, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b01100001; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01000010; c = 8'b00010100; // Expected: {'sum': 195, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01000010; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11100100; c = 8'b00110011; // Expected: {'sum': 66, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11100100; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b00011100; c = 8'b11100011; // Expected: {'sum': 148, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b00011100; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01110000; c = 8'b00001110; // Expected: {'sum': 254, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01110000; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10111100; c = 8'b10001001; // Expected: {'sum': 239, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10111100; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01110010; c = 8'b10111010; // Expected: {'sum': 73, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01110010; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00000111; c = 8'b11000011; // Expected: {'sum': 185, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00000111; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01001101; c = 8'b10101100; // Expected: {'sum': 56, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01001101; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10101100; c = 8'b11101010; // Expected: {'sum': 157, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10101100; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01001100; c = 8'b10110001; // Expected: {'sum': 86, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01001100; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10001010; c = 8'b00000111; // Expected: {'sum': 247, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10001010; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01000000; c = 8'b11010001; // Expected: {'sum': 210, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01000000; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11000100; c = 8'b10011011; // Expected: {'sum': 123, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11000100; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10111000; c = 8'b10000100; // Expected: {'sum': 136, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10111000; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01100110; c = 8'b01010100; // Expected: {'sum': 53, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01100110; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10011000; c = 8'b01010101; // Expected: {'sum': 54, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10011000; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10101001; c = 8'b10111101; // Expected: {'sum': 237, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10101001; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10100011; c = 8'b11110101; // Expected: {'sum': 144, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10100011; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00010111; c = 8'b10111100; // Expected: {'sum': 183, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00010111; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b01000110; c = 8'b00101111; // Expected: {'sum': 15, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b01000110; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10010110; c = 8'b10100111; // Expected: {'sum': 195, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10010110; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b00010001; c = 8'b11010011; // Expected: {'sum': 57, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b00010001; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01011100; c = 8'b11010110; // Expected: {'sum': 225, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01011100; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b11000111; c = 8'b10100111; // Expected: {'sum': 80, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b11000111; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11011100; c = 8'b00010010; // Expected: {'sum': 137, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11011100; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01100010; c = 8'b00001110; // Expected: {'sum': 15, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01100010; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00011010; c = 8'b01001010; // Expected: {'sum': 81, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00011010; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b10111000; c = 8'b10100111; // Expected: {'sum': 1, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b10111000; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b00110110; c = 8'b11111100; // Expected: {'sum': 165, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b00110110; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b01000110; c = 8'b00011000; // Expected: {'sum': 164, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b01000110; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01011000; c = 8'b11010000; // Expected: {'sum': 120, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01011000; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00110111; c = 8'b11100101; // Expected: {'sum': 35, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00110111; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10101110; c = 8'b00010011; // Expected: {'sum': 37, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10101110; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b00100000; c = 8'b10101110; // Expected: {'sum': 197, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b00100000; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00101100; c = 8'b00100100; // Expected: {'sum': 40, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00101100; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b01011111; c = 8'b01101101; // Expected: {'sum': 21, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b01011111; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10110100; c = 8'b00110001; // Expected: {'sum': 76, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10110100; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b00001000; c = 8'b11010111; // Expected: {'sum': 234, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b00001000; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11101110; c = 8'b01110001; // Expected: {'sum': 99, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11101110; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b10000100; c = 8'b01010010; // Expected: {'sum': 161, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b10000100; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b10110110; c = 8'b01001101; // Expected: {'sum': 102, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b10110110; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b01001100; c = 8'b10001110; // Expected: {'sum': 9, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b01001100; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00100110; c = 8'b00100100; // Expected: {'sum': 65, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00100110; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b10011011; c = 8'b11111000; // Expected: {'sum': 137, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b10011011; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10000110; c = 8'b11000110; // Expected: {'sum': 166, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10000110; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01010110; c = 8'b01000001; // Expected: {'sum': 11, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01010110; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01000000; c = 8'b10100001; // Expected: {'sum': 54, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01000000; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b11100111; c = 8'b01011000; // Expected: {'sum': 124, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b11100111; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10011010; c = 8'b10101100; // Expected: {'sum': 25, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10011010; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b10110101; c = 8'b11100111; // Expected: {'sum': 245, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b10110101; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10100001; c = 8'b01110001; // Expected: {'sum': 178, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10100001; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b11111011; c = 8'b00101100; // Expected: {'sum': 121, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b11111011; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b00011111; c = 8'b10101111; // Expected: {'sum': 139, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b00011111; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11101000; c = 8'b10111000; // Expected: {'sum': 16, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11101000; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00011000; c = 8'b11011101; // Expected: {'sum': 135, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00011000; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b10010001; c = 8'b00001000; // Expected: {'sum': 21, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b10010001; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10010101; c = 8'b00100010; // Expected: {'sum': 31, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10010101; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11000110; c = 8'b00110100; // Expected: {'sum': 237, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11000110; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b01101110; c = 8'b10101110; // Expected: {'sum': 39, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b01101110; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00001000; c = 8'b00001001; // Expected: {'sum': 205, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00001000; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b01010100; c = 8'b01011001; // Expected: {'sum': 212, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b01010100; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b00101001; c = 8'b10100111; // Expected: {'sum': 25, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b00101001; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10111011; c = 8'b00001100; // Expected: {'sum': 252, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10111011; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00010010; c = 8'b01010000; // Expected: {'sum': 39, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00010010; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b00110001; c = 8'b01110001; // Expected: {'sum': 163, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b00110001; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00111111; c = 8'b01110110; // Expected: {'sum': 73, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00111111; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00111010; c = 8'b11101110; // Expected: {'sum': 150, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00111010; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10111111; c = 8'b10110101; // Expected: {'sum': 238, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10111111; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10011011; c = 8'b11000001; // Expected: {'sum': 23, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10011011; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10100110; c = 8'b10100101; // Expected: {'sum': 73, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10100110; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10100110; c = 8'b01101010; // Expected: {'sum': 174, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10100110; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01011010; c = 8'b01010000; // Expected: {'sum': 169, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01011010; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10010010; c = 8'b01111011; // Expected: {'sum': 241, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10010010; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11100010; c = 8'b00110010; // Expected: {'sum': 152, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11100010; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00001011; c = 8'b01010100; // Expected: {'sum': 114, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00001011; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b00110101; c = 8'b00100011; // Expected: {'sum': 142, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b00110101; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b00110111; c = 8'b01111000; // Expected: {'sum': 192, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b00110111; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b11100000; c = 8'b11000000; // Expected: {'sum': 65, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b11100000; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b01011001; c = 8'b10111111; // Expected: {'sum': 209, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b01011001; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b00001100; c = 8'b00010110; // Expected: {'sum': 113, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b00001100; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01000111; c = 8'b01000110; // Expected: {'sum': 209, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01000111; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b00001100; c = 8'b11101110; // Expected: {'sum': 127, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b00001100; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01011000; c = 8'b10010010; // Expected: {'sum': 145, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01011000; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b01110110; c = 8'b00100000; // Expected: {'sum': 154, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b01110110; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01100010; c = 8'b10101000; // Expected: {'sum': 226, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01100010; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00010001; c = 8'b00110100; // Expected: {'sum': 173, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00010001; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b10001011; c = 8'b11101000; // Expected: {'sum': 205, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b10001011; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00100011; c = 8'b11100000; // Expected: {'sum': 224, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00100011; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11111111; c = 8'b11101010; // Expected: {'sum': 190, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11111111; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11011111; c = 8'b01111100; // Expected: {'sum': 222, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11011111; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b11010000; c = 8'b11111010; // Expected: {'sum': 239, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b11010000; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10110000; c = 8'b10010111; // Expected: {'sum': 84, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10110000; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11001111; c = 8'b00000001; // Expected: {'sum': 74, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11001111; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11101010; c = 8'b10111101; // Expected: {'sum': 115, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11101010; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b01110001; c = 8'b00101101; // Expected: {'sum': 107, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b01110001; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b01100100; c = 8'b00111100; // Expected: {'sum': 198, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b01100100; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11001100; c = 8'b10010011; // Expected: {'sum': 157, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11001100; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b01011111; c = 8'b00010001; // Expected: {'sum': 161, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b01011111; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11000000; c = 8'b00111011; // Expected: {'sum': 176, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11000000; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00010101; c = 8'b00101110; // Expected: {'sum': 59, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00010101; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00101001; c = 8'b11000000; // Expected: {'sum': 26, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00101001; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10101000; c = 8'b01001100; // Expected: {'sum': 129, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10101000; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01010000; c = 8'b11011100; // Expected: {'sum': 91, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01010000; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10000101; c = 8'b11111100; // Expected: {'sum': 34, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10000101; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10010010; c = 8'b00111000; // Expected: {'sum': 239, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10010010; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b01110110; c = 8'b01000110; // Expected: {'sum': 132, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b01110110; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b01010011; c = 8'b00011101; // Expected: {'sum': 164, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b01010011; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b00100111; c = 8'b01000110; // Expected: {'sum': 88, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b00100111; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10000011; c = 8'b00001110; // Expected: {'sum': 77, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10000011; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b00000011; c = 8'b01011111; // Expected: {'sum': 246, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b00000011; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00000100; c = 8'b00101010; // Expected: {'sum': 156, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00000100; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11111011; c = 8'b00101101; // Expected: {'sum': 78, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11111011; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b11110101; c = 8'b00111011; // Expected: {'sum': 175, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b11110101; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00101100; c = 8'b00000111; // Expected: {'sum': 77, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00101100; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b11010110; c = 8'b01110001; // Expected: {'sum': 87, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b11010110; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b11111001; c = 8'b11111000; // Expected: {'sum': 180, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b11111001; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b01001111; c = 8'b01101111; // Expected: {'sum': 237, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b01001111; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01101111; c = 8'b10000111; // Expected: {'sum': 84, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01101111; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b10000111; c = 8'b11011010; // Expected: {'sum': 179, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b10000111; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b00011001; c = 8'b01111101; // Expected: {'sum': 220, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b00011001; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10100110; c = 8'b00001111; // Expected: {'sum': 28, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10100110; c = 8'b00001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b11000001; c = 8'b01110101; // Expected: {'sum': 88, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b11000001; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01010011; c = 8'b11010000; // Expected: {'sum': 222, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01010011; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01111110; c = 8'b00000101; // Expected: {'sum': 38, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01111110; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b11101110; c = 8'b01101001; // Expected: {'sum': 74, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b11101110; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10010001; c = 8'b01010011; // Expected: {'sum': 144, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10010001; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10001101; c = 8'b10011010; // Expected: {'sum': 50, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10001101; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10010100; c = 8'b11011000; // Expected: {'sum': 144, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10010100; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11111011; c = 8'b00010011; // Expected: {'sum': 188, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11111011; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00011110; c = 8'b00001100; // Expected: {'sum': 50, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00011110; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b00111111; c = 8'b01000101; // Expected: {'sum': 104, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b00111111; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10111100; c = 8'b11010000; // Expected: {'sum': 191, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10111100; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b10010110; c = 8'b00001010; // Expected: {'sum': 46, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b10010110; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10100000; c = 8'b10110011; // Expected: {'sum': 9, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10100000; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10011101; c = 8'b00010111; // Expected: {'sum': 124, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10011101; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00111110; c = 8'b10101001; // Expected: {'sum': 11, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00111110; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b00001010; c = 8'b01100001; // Expected: {'sum': 183, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b00001010; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b00110110; c = 8'b01110111; // Expected: {'sum': 124, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b00110110; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b11000000; c = 8'b10010111; // Expected: {'sum': 196, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b11000000; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01011001; c = 8'b01110100; // Expected: {'sum': 195, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01011001; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b01101101; c = 8'b01101000; // Expected: {'sum': 211, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b01101101; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10100101; c = 8'b00001001; // Expected: {'sum': 110, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10100101; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b00011110; c = 8'b01101010; // Expected: {'sum': 67, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b00011110; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00110101; c = 8'b10011000; // Expected: {'sum': 79, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00110101; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b11101010; c = 8'b00111101; // Expected: {'sum': 139, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b11101010; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01110010; c = 8'b01111100; // Expected: {'sum': 203, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01110010; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01100000; c = 8'b10010100; // Expected: {'sum': 117, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01100000; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10111100; c = 8'b10001011; // Expected: {'sum': 49, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10111100; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b00101000; c = 8'b00111100; // Expected: {'sum': 70, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b00101000; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01100010; c = 8'b01011010; // Expected: {'sum': 151, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01100010; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10001101; c = 8'b00011010; // Expected: {'sum': 149, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10001101; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b00010101; c = 8'b10101101; // Expected: {'sum': 241, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b00010101; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10111000; c = 8'b01000000; // Expected: {'sum': 25, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10111000; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10100011; c = 8'b10001010; // Expected: {'sum': 145, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10100011; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00100010; c = 8'b00010011; // Expected: {'sum': 103, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00100010; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00011000; c = 8'b00111001; // Expected: {'sum': 92, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00011000; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10110010; c = 8'b11101001; // Expected: {'sum': 3, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10110010; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01010010; c = 8'b01000001; // Expected: {'sum': 164, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01010010; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10110110; c = 8'b11001001; // Expected: {'sum': 242, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10110110; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11100000; c = 8'b01000110; // Expected: {'sum': 128, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11100000; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b10111001; c = 8'b10100100; // Expected: {'sum': 228, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b10111001; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11111000; c = 8'b00000000; // Expected: {'sum': 203, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11111000; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b01111111; c = 8'b11110110; // Expected: {'sum': 86, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b01111111; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00000110; c = 8'b00110000; // Expected: {'sum': 80, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00000110; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00000110; c = 8'b01000010; // Expected: {'sum': 250, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00000110; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b00011000; c = 8'b11011110; // Expected: {'sum': 178, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b00011000; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00001000; c = 8'b10110000; // Expected: {'sum': 82, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00001000; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01000010; c = 8'b00110001; // Expected: {'sum': 1, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01000010; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11010000; c = 8'b01100110; // Expected: {'sum': 78, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11010000; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01111110; c = 8'b00100010; // Expected: {'sum': 250, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01111110; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00110111; c = 8'b00000110; // Expected: {'sum': 54, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00110111; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00111001; c = 8'b10010001; // Expected: {'sum': 35, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00111001; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b01101000; c = 8'b01000000; // Expected: {'sum': 73, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b01101000; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b11100000; c = 8'b11110111; // Expected: {'sum': 216, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b11100000; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10100000; c = 8'b11100001; // Expected: {'sum': 248, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10100000; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00101011; c = 8'b11101100; // Expected: {'sum': 131, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00101011; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11111001; c = 8'b00011100; // Expected: {'sum': 156, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11111001; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11110110; c = 8'b10001000; // Expected: {'sum': 5, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11110110; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01101001; c = 8'b00100100; // Expected: {'sum': 53, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01101001; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b00101110; c = 8'b10100101; // Expected: {'sum': 143, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b00101110; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10000000; c = 8'b10001001; // Expected: {'sum': 237, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10000000; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11101001; c = 8'b01101110; // Expected: {'sum': 21, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11101001; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10001000; c = 8'b10010111; // Expected: {'sum': 176, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10001000; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10010100; c = 8'b00101111; // Expected: {'sum': 79, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10010100; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00101111; c = 8'b10001111; // Expected: {'sum': 65, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00101111; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11000111; c = 8'b00011000; // Expected: {'sum': 117, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11000111; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11011001; c = 8'b01001101; // Expected: {'sum': 104, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11011001; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00010011; c = 8'b00001001; // Expected: {'sum': 127, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00010011; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11000101; c = 8'b00100100; // Expected: {'sum': 80, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11000101; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00011000; c = 8'b10010110; // Expected: {'sum': 151, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00011000; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b00011110; c = 8'b01001101; // Expected: {'sum': 21, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b00011110; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b11000000; c = 8'b00000001; // Expected: {'sum': 39, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b11000000; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1663,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b01110101; c = 8'b10010101; // Expected: {'sum': 251, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b01110101; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1664,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00101010; c = 8'b11110001; // Expected: {'sum': 128, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00101010; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1665,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11000000; c = 8'b10101111; // Expected: {'sum': 9, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11000000; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1666,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b00101101; c = 8'b00111101; // Expected: {'sum': 135, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b00101101; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1667,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00101001; c = 8'b00100000; // Expected: {'sum': 252, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00101001; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1668,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00010000; c = 8'b11111111; // Expected: {'sum': 89, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00010000; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1669,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00001100; c = 8'b00111001; // Expected: {'sum': 100, 'carry': 25}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00001100; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1670,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b10110010; c = 8'b01000111; // Expected: {'sum': 18, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b10110010; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1671,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b11110010; c = 8'b01101101; // Expected: {'sum': 34, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b11110010; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1672,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b11011110; c = 8'b10110100; // Expected: {'sum': 240, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b11011110; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1673,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10010111; c = 8'b11101001; // Expected: {'sum': 224, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10010111; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1674,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10011111; c = 8'b11101010; // Expected: {'sum': 104, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10011111; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1675,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b11100000; c = 8'b00010111; // Expected: {'sum': 21, 'carry': 226}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b11100000; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1676,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b11110011; c = 8'b00011000; // Expected: {'sum': 39, 'carry': 216}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b11110011; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1677,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00100110; c = 8'b00001101; // Expected: {'sum': 76, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00100110; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1678,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b11010010; c = 8'b00111100; // Expected: {'sum': 114, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b11010010; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1679,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b01111001; c = 8'b11000000; // Expected: {'sum': 12, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b01111001; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1680,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01000100; c = 8'b00011101; // Expected: {'sum': 214, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01000100; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1681,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10100110; c = 8'b01001000; // Expected: {'sum': 253, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10100110; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1682,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11000001; c = 8'b00010011; // Expected: {'sum': 120, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11000001; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1683,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11100110; c = 8'b11010000; // Expected: {'sum': 138, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11100110; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1684,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b01110110; c = 8'b01011010; // Expected: {'sum': 166, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b01110110; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1685,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11011110; c = 8'b00110101; // Expected: {'sum': 15, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11011110; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1686,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b11110010; c = 8'b10001111; // Expected: {'sum': 97, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b11110010; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1687,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10101111; c = 8'b00110111; // Expected: {'sum': 184, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10101111; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1688,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11001110; c = 8'b10010101; // Expected: {'sum': 22, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11001110; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1689,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01100111; c = 8'b11011011; // Expected: {'sum': 81, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01100111; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1690,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00011111; c = 8'b00101100; // Expected: {'sum': 68, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00011111; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1691,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10000010; c = 8'b00001011; // Expected: {'sum': 52, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10000010; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1692,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01001001; c = 8'b00000101; // Expected: {'sum': 122, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01001001; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1693,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10111000; c = 8'b11001000; // Expected: {'sum': 156, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10111000; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1694,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b11110100; c = 8'b10000100; // Expected: {'sum': 185, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b11110100; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1695,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b10001100; c = 8'b00000101; // Expected: {'sum': 252, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b10001100; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1696,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b01001011; c = 8'b11000010; // Expected: {'sum': 138, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b01001011; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1697,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10111001; c = 8'b00010101; // Expected: {'sum': 186, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10111001; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1698,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b11111001; c = 8'b11111011; // Expected: {'sum': 233, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b11111001; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1699,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00001001; c = 8'b00111101; // Expected: {'sum': 81, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00001001; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1700,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01101101; c = 8'b01100000; // Expected: {'sum': 205, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01101101; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1701,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b11011111; c = 8'b11001000; // Expected: {'sum': 160, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b11011111; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1702,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01100010; c = 8'b01100011; // Expected: {'sum': 61, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01100010; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1703,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b11000001; c = 8'b11010110; // Expected: {'sum': 249, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b11000001; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1704,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b11000101; c = 8'b00100010; // Expected: {'sum': 136, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b11000101; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1705,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00011111; c = 8'b01111011; // Expected: {'sum': 21, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00011111; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1706,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00111011; c = 8'b10101010; // Expected: {'sum': 65, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00111011; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1707,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b11111001; c = 8'b01110000; // Expected: {'sum': 43, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b11111001; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1708,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00010011; c = 8'b00001110; // Expected: {'sum': 117, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00010011; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1709,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01100001; c = 8'b00111010; // Expected: {'sum': 203, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01100001; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1710,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b10011100; c = 8'b00000010; // Expected: {'sum': 177, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b10011100; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1711,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b11100100; c = 8'b11000110; // Expected: {'sum': 251, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b11100100; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1712,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01111001; c = 8'b10100010; // Expected: {'sum': 160, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01111001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1713,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01100111; c = 8'b10111001; // Expected: {'sum': 138, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01100111; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1714,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11000101; c = 8'b11100001; // Expected: {'sum': 168, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11000101; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1715,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00001001; c = 8'b10100110; // Expected: {'sum': 156, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00001001; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1716,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10101011; c = 8'b00011000; // Expected: {'sum': 228, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10101011; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1717,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00000001; c = 8'b11001010; // Expected: {'sum': 90, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00000001; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1718,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01110001; c = 8'b10100111; // Expected: {'sum': 138, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01110001; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1719,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11101101; c = 8'b01110001; // Expected: {'sum': 225, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11101101; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1720,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01010110; c = 8'b10001101; // Expected: {'sum': 113, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01010110; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1721,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10011110; c = 8'b11111001; // Expected: {'sum': 107, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10011110; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1722,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01110101; c = 8'b00001101; // Expected: {'sum': 80, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01110101; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1723,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11011111; c = 8'b10011110; // Expected: {'sum': 150, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11011111; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1724,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11001111; c = 8'b00000100; // Expected: {'sum': 79, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11001111; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1725,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10000101; c = 8'b10010100; // Expected: {'sum': 52, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10000101; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1726,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10110010; c = 8'b01101000; // Expected: {'sum': 9, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10110010; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1727,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b00101010; c = 8'b10110110; // Expected: {'sum': 127, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b00101010; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1728,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11111000; c = 8'b10110000; // Expected: {'sum': 144, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11111000; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1729,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00011011; c = 8'b11010011; // Expected: {'sum': 114, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00011011; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1730,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01010110; c = 8'b10000110; // Expected: {'sum': 108, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01010110; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1731,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11101010; c = 8'b00101011; // Expected: {'sum': 3, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11101010; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1732,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11000011; c = 8'b11100011; // Expected: {'sum': 98, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11000011; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1733,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10001110; c = 8'b00111000; // Expected: {'sum': 247, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10001110; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1734,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b00001011; c = 8'b00101110; // Expected: {'sum': 154, 'carry': 47}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b00001011; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1735,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00101010; c = 8'b10011111; // Expected: {'sum': 54, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00101010; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1736,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b01111010; c = 8'b10000011; // Expected: {'sum': 3, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b01111010; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1737,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01000001; c = 8'b10011011; // Expected: {'sum': 2, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01000001; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1738,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b10111000; c = 8'b01010111; // Expected: {'sum': 234, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b10111000; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1739,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11110000; c = 8'b11110001; // Expected: {'sum': 84, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11110000; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1740,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10100101; c = 8'b01000011; // Expected: {'sum': 252, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10100101; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1741,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00111100; c = 8'b11100100; // Expected: {'sum': 43, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00111100; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1742,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10011110; c = 8'b01011100; // Expected: {'sum': 118, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10011110; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1743,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11011010; c = 8'b00011111; // Expected: {'sum': 240, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11011010; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1744,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00011101; c = 8'b00010000; // Expected: {'sum': 162, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00011101; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1745,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b11111010; c = 8'b00110001; // Expected: {'sum': 116, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b11111010; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1746,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01101010; c = 8'b00001001; // Expected: {'sum': 75, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01101010; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1747,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b11100001; c = 8'b10001001; // Expected: {'sum': 60, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b11100001; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1748,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b10011111; c = 8'b11010110; // Expected: {'sum': 223, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b10011111; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1749,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110010; c = 8'b11100110; // Expected: {'sum': 246, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110010; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1750,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01000010; c = 8'b01000000; // Expected: {'sum': 22, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01000010; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1751,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b10111000; c = 8'b11010101; // Expected: {'sum': 69, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b10111000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1752,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11101100; c = 8'b01011001; // Expected: {'sum': 228, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11101100; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1753,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b11111001; c = 8'b00001000; // Expected: {'sum': 48, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b11111001; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1754,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11110110; c = 8'b01111001; // Expected: {'sum': 235, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11110110; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1755,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11000001; c = 8'b01000111; // Expected: {'sum': 52, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11000001; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1756,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00001101; c = 8'b10100011; // Expected: {'sum': 20, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00001101; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1757,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01101001; c = 8'b00101010; // Expected: {'sum': 1, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01101001; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1758,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01010010; c = 8'b01001010; // Expected: {'sum': 33, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01010010; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1759,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01111100; c = 8'b11010001; // Expected: {'sum': 69, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01111100; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1760,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10100001; c = 8'b01001111; // Expected: {'sum': 50, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10100001; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1761,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00010000; c = 8'b01111000; // Expected: {'sum': 191, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00010000; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1762,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b11110011; c = 8'b00000001; // Expected: {'sum': 68, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b11110011; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1763,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b01000001; c = 8'b01011010; // Expected: {'sum': 36, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b01000001; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1764,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11001001; c = 8'b01011011; // Expected: {'sum': 46, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11001001; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1765,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10010100; c = 8'b10010011; // Expected: {'sum': 192, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10010100; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1766,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11111010; c = 8'b01111000; // Expected: {'sum': 51, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11111010; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1767,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b00111011; c = 8'b00011101; // Expected: {'sum': 145, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b00111011; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1768,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11010011; c = 8'b01100001; // Expected: {'sum': 242, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11010011; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1769,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10110101; c = 8'b10011111; // Expected: {'sum': 230, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10110101; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1770,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b00011110; c = 8'b00000000; // Expected: {'sum': 180, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b00011110; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1771,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01111100; c = 8'b00010110; // Expected: {'sum': 145, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01111100; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1772,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b00111101; c = 8'b10010001; // Expected: {'sum': 151, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b00111101; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1773,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00010000; c = 8'b01111010; // Expected: {'sum': 88, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00010000; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1774,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00101111; c = 8'b11101001; // Expected: {'sum': 33, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00101111; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1775,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b00001010; c = 8'b10100111; // Expected: {'sum': 223, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b00001010; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1776,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10000000; c = 8'b01011110; // Expected: {'sum': 130, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10000000; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1777,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10001011; c = 8'b11010000; // Expected: {'sum': 244, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10001011; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1778,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01101111; c = 8'b11001001; // Expected: {'sum': 253, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01101111; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1779,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10110101; c = 8'b01001111; // Expected: {'sum': 92, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10110101; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1780,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b11010011; c = 8'b10101000; // Expected: {'sum': 31, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b11010011; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1781,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01111000; c = 8'b10000000; // Expected: {'sum': 236, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01111000; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1782,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00011011; c = 8'b10001111; // Expected: {'sum': 160, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00011011; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1783,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b00011110; c = 8'b10110110; // Expected: {'sum': 222, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b00011110; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1784,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b11011111; c = 8'b01001001; // Expected: {'sum': 233, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b11011111; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1785,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00001110; c = 8'b10110001; // Expected: {'sum': 242, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00001110; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1786,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b01011000; c = 8'b00110011; // Expected: {'sum': 228, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b01011000; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1787,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10010000; c = 8'b01011101; // Expected: {'sum': 117, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10010000; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1788,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01001101; c = 8'b00011010; // Expected: {'sum': 192, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01001101; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1789,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01000000; c = 8'b11011011; // Expected: {'sum': 105, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01000000; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1790,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11100011; c = 8'b10110000; // Expected: {'sum': 127, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11100011; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1791,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01000001; c = 8'b11101000; // Expected: {'sum': 10, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01000001; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1792,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10100000; c = 8'b00101010; // Expected: {'sum': 130, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10100000; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1793,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10001111; c = 8'b01111100; // Expected: {'sum': 97, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10001111; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1794,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01011000; c = 8'b00101111; // Expected: {'sum': 83, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01011000; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1795,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b00101100; c = 8'b10001010; // Expected: {'sum': 71, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b00101100; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1796,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00110110; c = 8'b00010010; // Expected: {'sum': 212, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00110110; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1797,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00101101; c = 8'b01110101; // Expected: {'sum': 206, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00101101; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1798,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01110011; c = 8'b10110111; // Expected: {'sum': 111, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01110011; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1799,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b11011000; c = 8'b00000010; // Expected: {'sum': 116, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b11011000; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1800,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b10111100; c = 8'b01100001; // Expected: {'sum': 193, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b10111100; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1801,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b00000100; c = 8'b11110111; // Expected: {'sum': 147, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b00000100; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1802,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10010001; c = 8'b00010010; // Expected: {'sum': 163, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10010001; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1803,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11111010; c = 8'b01111111; // Expected: {'sum': 96, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11111010; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1804,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00000001; c = 8'b00000000; // Expected: {'sum': 63, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00000001; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1805,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11111011; c = 8'b11111101; // Expected: {'sum': 65, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11111011; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1806,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00111111; c = 8'b10000000; // Expected: {'sum': 111, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00111111; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1807,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00101010; c = 8'b00110010; // Expected: {'sum': 205, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00101010; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1808,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00100100; c = 8'b01000011; // Expected: {'sum': 85, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00100100; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1809,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b01111010; c = 8'b01110111; // Expected: {'sum': 22, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b01111010; c = 8'b01110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1810,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b01010011; c = 8'b10010010; // Expected: {'sum': 30, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b01010011; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1811,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11101010; c = 8'b10001101; // Expected: {'sum': 100, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11101010; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1812,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b10100000; c = 8'b10001100; // Expected: {'sum': 94, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b10100000; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1813,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b01000000; c = 8'b01010100; // Expected: {'sum': 150, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b01000000; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1814,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01010001; c = 8'b11010010; // Expected: {'sum': 58, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01010001; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1815,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11001110; c = 8'b11100100; // Expected: {'sum': 31, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11001110; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1816,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00011011; c = 8'b11110011; // Expected: {'sum': 29, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00011011; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1817,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b00101111; c = 8'b00111100; // Expected: {'sum': 2, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b00101111; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1818,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b11111111; c = 8'b01000100; // Expected: {'sum': 169, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b11111111; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1819,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11011111; c = 8'b11011110; // Expected: {'sum': 34, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11011111; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1820,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b10110100; c = 8'b00100011; // Expected: {'sum': 88, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b10110100; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1821,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b01100000; c = 8'b00000010; // Expected: {'sum': 189, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b01100000; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1822,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10111010; c = 8'b11000101; // Expected: {'sum': 178, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10111010; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1823,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10111110; c = 8'b00001001; // Expected: {'sum': 44, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10111110; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1824,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b11011100; c = 8'b00111001; // Expected: {'sum': 212, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b11011100; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1825,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b11000000; c = 8'b10000011; // Expected: {'sum': 14, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b11000000; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1826,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00110011; c = 8'b00101011; // Expected: {'sum': 40, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00110011; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1827,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11100110; c = 8'b11111111; // Expected: {'sum': 89, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11100110; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1828,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01001100; c = 8'b10100000; // Expected: {'sum': 8, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01001100; c = 8'b10100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1829,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10001011; c = 8'b01010000; // Expected: {'sum': 45, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10001011; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1830,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10111000; c = 8'b10010010; // Expected: {'sum': 137, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10111000; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1831,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01011011; c = 8'b01111111; // Expected: {'sum': 46, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01011011; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1832,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b10011100; c = 8'b11110000; // Expected: {'sum': 208, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b10011100; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1833,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01001100; c = 8'b00001010; // Expected: {'sum': 231, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01001100; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1834,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b10000100; c = 8'b00101110; // Expected: {'sum': 17, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b10000100; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1835,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b00101110; c = 8'b01011011; // Expected: {'sum': 211, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b00101110; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1836,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11101101; c = 8'b00101000; // Expected: {'sum': 167, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11101101; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1837,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01101110; c = 8'b01011011; // Expected: {'sum': 107, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01101110; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1838,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10000100; c = 8'b10010101; // Expected: {'sum': 97, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10000100; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1839,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b11010000; c = 8'b10101001; // Expected: {'sum': 108, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b11010000; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1840,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11011000; c = 8'b01000011; // Expected: {'sum': 22, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11011000; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1841,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10101110; c = 8'b00101001; // Expected: {'sum': 71, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10101110; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1842,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b01101001; c = 8'b01011011; // Expected: {'sum': 13, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b01101001; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1843,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01010101; c = 8'b11001111; // Expected: {'sum': 169, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01010101; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1844,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10111101; c = 8'b00111110; // Expected: {'sum': 0, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10111101; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1845,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10111000; c = 8'b00010011; // Expected: {'sum': 231, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10111000; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1846,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01011110; c = 8'b01111100; // Expected: {'sum': 139, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01011110; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1847,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11000111; c = 8'b00111011; // Expected: {'sum': 100, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11000111; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1848,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b00011000; c = 8'b10100111; // Expected: {'sum': 244, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b00011000; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1849,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b10111111; c = 8'b00100010; // Expected: {'sum': 239, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b10111111; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1850,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00100100; c = 8'b01001010; // Expected: {'sum': 15, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00100100; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1851,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b11111000; c = 8'b01010100; // Expected: {'sum': 81, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b11111000; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1852,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01101101; c = 8'b00110011; // Expected: {'sum': 34, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01101101; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1853,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b11010101; c = 8'b11101001; // Expected: {'sum': 155, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b11010101; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1854,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00100111; c = 8'b10110100; // Expected: {'sum': 45, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00100111; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1855,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11111101; c = 8'b10100001; // Expected: {'sum': 196, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11111101; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1856,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b00111101; c = 8'b01000110; // Expected: {'sum': 48, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b00111101; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1857,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00100001; c = 8'b10101101; // Expected: {'sum': 33, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00100001; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1858,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00110010; c = 8'b11110110; // Expected: {'sum': 153, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00110010; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1859,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11010010; c = 8'b10101010; // Expected: {'sum': 210, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11010010; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1860,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b10111001; c = 8'b00111101; // Expected: {'sum': 27, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b10111001; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1861,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01101011; c = 8'b01110110; // Expected: {'sum': 29, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01101011; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1862,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b01011010; c = 8'b11100010; // Expected: {'sum': 131, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b01011010; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1863,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11011010; c = 8'b10011111; // Expected: {'sum': 72, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11011010; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1864,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00111001; c = 8'b00111010; // Expected: {'sum': 137, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00111001; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1865,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01101101; c = 8'b00010110; // Expected: {'sum': 38, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01101101; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1866,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11010101; c = 8'b01000110; // Expected: {'sum': 3, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11010101; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1867,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01000111; c = 8'b01010010; // Expected: {'sum': 49, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01000111; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1868,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11110101; c = 8'b11100010; // Expected: {'sum': 3, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11110101; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1869,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b01011111; c = 8'b00110001; // Expected: {'sum': 221, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b01011111; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1870,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b11010111; c = 8'b11001100; // Expected: {'sum': 20, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b11010111; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1871,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01100011; c = 8'b00001010; // Expected: {'sum': 177, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01100011; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1872,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11101100; c = 8'b01100101; // Expected: {'sum': 45, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11101100; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1873,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01000001; c = 8'b00111010; // Expected: {'sum': 71, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01000001; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1874,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11000011; c = 8'b10111000; // Expected: {'sum': 208, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11000011; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1875,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10010000; c = 8'b00011010; // Expected: {'sum': 198, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10010000; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1876,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b01000001; c = 8'b11100101; // Expected: {'sum': 153, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b01000001; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1877,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b01000111; c = 8'b10010000; // Expected: {'sum': 205, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b01000111; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1878,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10110111; c = 8'b01011110; // Expected: {'sum': 18, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10110111; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1879,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01111000; c = 8'b11110011; // Expected: {'sum': 184, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01111000; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1880,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b01011001; c = 8'b10100100; // Expected: {'sum': 182, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b01011001; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1881,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b10011111; c = 8'b01010000; // Expected: {'sum': 28, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b10011111; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1882,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00001010; c = 8'b01101010; // Expected: {'sum': 5, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00001010; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1883,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b11010101; c = 8'b01001001; // Expected: {'sum': 97, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b11010101; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1884,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01101111; c = 8'b00011111; // Expected: {'sum': 52, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01101111; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1885,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b11101000; c = 8'b10000010; // Expected: {'sum': 118, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b11101000; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1886,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b01100001; c = 8'b01001101; // Expected: {'sum': 125, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b01100001; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1887,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11100111; c = 8'b01101100; // Expected: {'sum': 156, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11100111; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1888,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b11001001; c = 8'b01101001; // Expected: {'sum': 255, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b11001001; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1889,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10000010; c = 8'b10001111; // Expected: {'sum': 55, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10000010; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1890,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b01010110; c = 8'b00100010; // Expected: {'sum': 113, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b01010110; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1891,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b01010001; c = 8'b00000000; // Expected: {'sum': 166, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b01010001; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1892,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10011110; c = 8'b00100010; // Expected: {'sum': 225, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10011110; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1893,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b00110010; c = 8'b11111001; // Expected: {'sum': 33, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b00110010; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1894,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11010101; c = 8'b11100011; // Expected: {'sum': 62, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11010101; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1895,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b01111001; c = 8'b00011000; // Expected: {'sum': 19, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b01111001; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1896,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11110001; c = 8'b10100001; // Expected: {'sum': 250, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11110001; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1897,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b11001101; c = 8'b11110011; // Expected: {'sum': 58, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b11001101; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1898,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b11110101; c = 8'b01101011; // Expected: {'sum': 64, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b11110101; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1899,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b01001110; c = 8'b01001001; // Expected: {'sum': 28, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b01001110; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1900,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00101011; c = 8'b10110110; // Expected: {'sum': 108, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00101011; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1901,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b00011000; c = 8'b01000111; // Expected: {'sum': 97, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b00011000; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1902,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01010011; c = 8'b01110100; // Expected: {'sum': 139, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01010011; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1903,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10101000; c = 8'b11011110; // Expected: {'sum': 244, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10101000; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1904,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b00010111; c = 8'b10111101; // Expected: {'sum': 184, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b00010111; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1905,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11001101; c = 8'b10011100; // Expected: {'sum': 195, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11001101; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1906,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b01000010; c = 8'b10000001; // Expected: {'sum': 207, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b01000010; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1907,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01000011; c = 8'b11001000; // Expected: {'sum': 73, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01000011; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1908,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00010100; c = 8'b11101110; // Expected: {'sum': 223, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00010100; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1909,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01100001; c = 8'b11001001; // Expected: {'sum': 196, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01100001; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1910,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01101011; c = 8'b01000100; // Expected: {'sum': 5, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01101011; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1911,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00011111; c = 8'b00011100; // Expected: {'sum': 199, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00011111; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1912,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00000111; c = 8'b01100101; // Expected: {'sum': 211, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00000111; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1913,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10000000; c = 8'b01100101; // Expected: {'sum': 116, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10000000; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1914,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10110101; c = 8'b01100001; // Expected: {'sum': 164, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10110101; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1915,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00010000; c = 8'b01001111; // Expected: {'sum': 238, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00010000; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1916,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11101101; c = 8'b01011001; // Expected: {'sum': 142, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11101101; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1917,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01001111; c = 8'b10010101; // Expected: {'sum': 63, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01001111; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1918,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00110100; c = 8'b10101011; // Expected: {'sum': 20, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00110100; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1919,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10110101; c = 8'b01010101; // Expected: {'sum': 90, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10110101; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1920,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11110000; c = 8'b01011001; // Expected: {'sum': 212, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11110000; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1921,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b10110000; c = 8'b01011011; // Expected: {'sum': 121, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b10110000; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1922,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b00010011; c = 8'b11001011; // Expected: {'sum': 238, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b00010011; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1923,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b00000100; c = 8'b01111011; // Expected: {'sum': 180, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b00000100; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1924,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11010100; c = 8'b10010000; // Expected: {'sum': 204, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11010100; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1925,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01000010; c = 8'b00111011; // Expected: {'sum': 26, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01000010; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1926,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01101110; c = 8'b01101001; // Expected: {'sum': 62, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01101110; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1927,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b10110010; c = 8'b00001111; // Expected: {'sum': 159, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b10110010; c = 8'b00001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1928,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b01100001; c = 8'b01110101; // Expected: {'sum': 248, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b01100001; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1929,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b00110110; c = 8'b01000000; // Expected: {'sum': 206, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b00110110; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1930,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b10011101; c = 8'b00011111; // Expected: {'sum': 84, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b10011101; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1931,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b11111001; c = 8'b11010110; // Expected: {'sum': 83, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b11111001; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1932,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b10011100; c = 8'b01011101; // Expected: {'sum': 230, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b10011100; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1933,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b10010001; c = 8'b10111010; // Expected: {'sum': 224, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b10010001; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1934,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00110111; c = 8'b01010110; // Expected: {'sum': 159, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00110111; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1935,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b11110001; c = 8'b00011001; // Expected: {'sum': 234, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b11110001; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1936,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10000100; c = 8'b11011001; // Expected: {'sum': 177, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10000100; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1937,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b10110101; c = 8'b01100001; // Expected: {'sum': 242, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b10110101; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1938,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11110111; c = 8'b00001011; // Expected: {'sum': 137, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11110111; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1939,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10011111; c = 8'b00001101; // Expected: {'sum': 59, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10011111; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1940,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11111011; c = 8'b01101001; // Expected: {'sum': 201, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11111011; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1941,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b11111010; c = 8'b00011010; // Expected: {'sum': 104, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b11111010; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1942,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b01000100; c = 8'b01101110; // Expected: {'sum': 164, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b01000100; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1943,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b10011110; c = 8'b10010111; // Expected: {'sum': 127, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b10011110; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1944,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01100111; c = 8'b11010111; // Expected: {'sum': 128, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01100111; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1945,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11101110; c = 8'b11001011; // Expected: {'sum': 49, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11101110; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1946,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10100000; c = 8'b10110101; // Expected: {'sum': 72, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10100000; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1947,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11111011; c = 8'b11010000; // Expected: {'sum': 128, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11111011; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1948,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01010101; c = 8'b01010000; // Expected: {'sum': 188, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01010101; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1949,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00011110; c = 8'b10000110; // Expected: {'sum': 168, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00011110; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1950,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01111100; c = 8'b01001100; // Expected: {'sum': 160, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01111100; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1951,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10101010; c = 8'b10001110; // Expected: {'sum': 246, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10101010; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1952,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b11100111; c = 8'b01111010; // Expected: {'sum': 9, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b11100111; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1953,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00011001; c = 8'b10000000; // Expected: {'sum': 146, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00011001; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1954,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b10100110; c = 8'b00100100; // Expected: {'sum': 50, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b10100110; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1955,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10100010; c = 8'b01101000; // Expected: {'sum': 227, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10100010; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1956,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00001000; c = 8'b01111110; // Expected: {'sum': 215, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00001000; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1957,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b11010100; c = 8'b11100101; // Expected: {'sum': 193, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b11010100; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1958,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01001000; c = 8'b10111011; // Expected: {'sum': 152, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01001000; c = 8'b10111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1959,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00001001; c = 8'b10000001; // Expected: {'sum': 100, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00001001; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1960,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00001100; c = 8'b10111001; // Expected: {'sum': 217, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00001100; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1961,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01100001; c = 8'b11010101; // Expected: {'sum': 52, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01100001; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1962,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b11101110; c = 8'b00001000; // Expected: {'sum': 25, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b11101110; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1963,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00110101; c = 8'b11100001; // Expected: {'sum': 171, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00110101; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1964,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01000001; c = 8'b10011110; // Expected: {'sum': 188, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01000001; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1965,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01111000; c = 8'b11010101; // Expected: {'sum': 100, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01111000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1966,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01000110; c = 8'b01111111; // Expected: {'sum': 45, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01000110; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1967,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b10100010; c = 8'b00110010; // Expected: {'sum': 102, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b10100010; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1968,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b00001010; c = 8'b11011010; // Expected: {'sum': 239, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b00001010; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1969,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b10111011; c = 8'b10111001; // Expected: {'sum': 40, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b10111011; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1970,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b00011100; c = 8'b11111110; // Expected: {'sum': 164, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b00011100; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1971,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10100101; c = 8'b01100100; // Expected: {'sum': 236, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10100101; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1972,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b01000000; c = 8'b10001110; // Expected: {'sum': 222, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b01000000; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1973,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01101111; c = 8'b10110000; // Expected: {'sum': 155, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01101111; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1974,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10010000; c = 8'b00100010; // Expected: {'sum': 133, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10010000; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1975,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01100011; c = 8'b10110111; // Expected: {'sum': 70, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01100011; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1976,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01001110; c = 8'b11110001; // Expected: {'sum': 220, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01001110; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1977,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10100100; c = 8'b01000001; // Expected: {'sum': 225, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10100100; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1978,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10011011; c = 8'b00111100; // Expected: {'sum': 125, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10011011; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1979,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11000011; c = 8'b00111100; // Expected: {'sum': 110, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11000011; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1980,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01110000; c = 8'b00110000; // Expected: {'sum': 205, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01110000; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1981,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00101000; c = 8'b10110101; // Expected: {'sum': 27, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00101000; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1982,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01000111; c = 8'b00111000; // Expected: {'sum': 247, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01000111; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1983,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00100011; c = 8'b00111111; // Expected: {'sum': 11, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00100011; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1984,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01001010; c = 8'b10100101; // Expected: {'sum': 139, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01001010; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1985,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11100101; c = 8'b00001100; // Expected: {'sum': 188, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11100101; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1986,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b00100110; c = 8'b10100111; // Expected: {'sum': 94, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b00100110; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1987,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01100110; c = 8'b10101011; // Expected: {'sum': 110, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01100110; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1988,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00110101; c = 8'b00100101; // Expected: {'sum': 181, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00110101; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1989,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11111001; c = 8'b00001110; // Expected: {'sum': 169, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11111001; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1990,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b01111000; c = 8'b00111011; // Expected: {'sum': 145, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b01111000; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1991,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01000011; c = 8'b11110111; // Expected: {'sum': 12, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01000011; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1992,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10101100; c = 8'b11111111; // Expected: {'sum': 238, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10101100; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1993,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10101111; c = 8'b10110110; // Expected: {'sum': 151, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10101111; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1994,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11000010; c = 8'b00111001; // Expected: {'sum': 142, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11000010; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1995,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10001101; c = 8'b10111011; // Expected: {'sum': 221, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10001101; c = 8'b10111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1996,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11001110; c = 8'b00101101; // Expected: {'sum': 143, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11001110; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1997,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10110000; c = 8'b10110100; // Expected: {'sum': 252, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10110000; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1998,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11010101; c = 8'b01011000; // Expected: {'sum': 184, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11010101; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1999,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11100011; c = 8'b10110100; // Expected: {'sum': 38, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11100011; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2000,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10110001; c = 8'b10100010; // Expected: {'sum': 41, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10110001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2001,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01111100; c = 8'b11110000; // Expected: {'sum': 212, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01111100; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2002,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00000101; c = 8'b00110010; // Expected: {'sum': 137, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00000101; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2003,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00010001; c = 8'b00111011; // Expected: {'sum': 68, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00010001; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2004,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01101101; c = 8'b11000011; // Expected: {'sum': 146, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01101101; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2005,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b01110000; c = 8'b01100001; // Expected: {'sum': 20, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b01110000; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2006,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00001001; c = 8'b11010000; // Expected: {'sum': 187, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00001001; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2007,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11100111; c = 8'b11110110; // Expected: {'sum': 140, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11100111; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2008,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00110100; c = 8'b01000011; // Expected: {'sum': 220, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00110100; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2009,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01101000; c = 8'b11000001; // Expected: {'sum': 60, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01101000; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2010,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11110110; c = 8'b01000111; // Expected: {'sum': 224, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11110110; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2011,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b01111011; c = 8'b00010110; // Expected: {'sum': 222, 'carry': 51}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b01111011; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2012,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11000110; c = 8'b10010100; // Expected: {'sum': 126, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11000110; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2013,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10010011; c = 8'b01100101; // Expected: {'sum': 27, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10010011; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2014,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b01011111; c = 8'b10110110; // Expected: {'sum': 120, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b01011111; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2015,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01000110; c = 8'b00001100; // Expected: {'sum': 253, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01000110; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2016,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01100111; c = 8'b00001100; // Expected: {'sum': 16, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01100111; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2017,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00001010; c = 8'b10110001; // Expected: {'sum': 185, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00001010; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2018,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11100000; c = 8'b00111110; // Expected: {'sum': 83, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11100000; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2019,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10111101; c = 8'b01010000; // Expected: {'sum': 131, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10111101; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2020,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00001110; c = 8'b11011100; // Expected: {'sum': 5, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00001110; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2021,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11001011; c = 8'b11011000; // Expected: {'sum': 42, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11001011; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2022,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b10010111; c = 8'b01101101; // Expected: {'sum': 155, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b10010111; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2023,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11111001; c = 8'b11011011; // Expected: {'sum': 72, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11111001; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2024,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00110111; c = 8'b01111010; // Expected: {'sum': 131, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00110111; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2025,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01000111; c = 8'b01101111; // Expected: {'sum': 243, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01000111; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2026,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10110101; c = 8'b00011010; // Expected: {'sum': 193, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10110101; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2027,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b00100111; c = 8'b00000111; // Expected: {'sum': 173, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b00100111; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2028,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b01000100; c = 8'b10111010; // Expected: {'sum': 240, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b01000100; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2029,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b11111001; c = 8'b10101100; // Expected: {'sum': 82, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b11111001; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2030,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00111101; c = 8'b11000101; // Expected: {'sum': 230, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00111101; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2031,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b00000101; c = 8'b11111110; // Expected: {'sum': 95, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b00000101; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2032,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b01000000; c = 8'b11111111; // Expected: {'sum': 203, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b01000000; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2033,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10101110; c = 8'b00110101; // Expected: {'sum': 63, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10101110; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2034,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11001110; c = 8'b01101010; // Expected: {'sum': 37, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11001110; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2035,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b11100011; c = 8'b11010001; // Expected: {'sum': 173, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b11100011; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2036,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00010110; c = 8'b10011111; // Expected: {'sum': 120, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00010110; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2037,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b00001000; c = 8'b11100111; // Expected: {'sum': 123, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b00001000; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2038,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00000000; c = 8'b01010000; // Expected: {'sum': 128, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00000000; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2039,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01111001; c = 8'b01000001; // Expected: {'sum': 67, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01111001; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2040,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00010100; c = 8'b01101110; // Expected: {'sum': 20, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00010100; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2041,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11110110; c = 8'b10111010; // Expected: {'sum': 21, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11110110; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2042,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11010011; c = 8'b00100101; // Expected: {'sum': 15, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11010011; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2043,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b11010111; c = 8'b11010000; // Expected: {'sum': 188, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b11010111; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2044,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b01100011; c = 8'b11110101; // Expected: {'sum': 80, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b01100011; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2045,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10111110; c = 8'b00000010; // Expected: {'sum': 215, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10111110; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2046,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b01110111; c = 8'b01010010; // Expected: {'sum': 220, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b01110111; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2047,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00111001; c = 8'b00001110; // Expected: {'sum': 154, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00111001; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2048,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b11001110; c = 8'b10101100; // Expected: {'sum': 206, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b11001110; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2049,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00010000; c = 8'b01101011; // Expected: {'sum': 90, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00010000; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2050,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00101111; c = 8'b00100110; // Expected: {'sum': 44, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00101111; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2051,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b11111100; c = 8'b01101110; // Expected: {'sum': 87, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b11111100; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2052,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b10111111; c = 8'b10001010; // Expected: {'sum': 190, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b10111111; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2053,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10001111; c = 8'b11100000; // Expected: {'sum': 70, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10001111; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2054,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b01101110; c = 8'b10011111; // Expected: {'sum': 136, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b01101110; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2055,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10000010; c = 8'b11000110; // Expected: {'sum': 3, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10000010; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2056,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b11000011; c = 8'b01110000; // Expected: {'sum': 84, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b11000011; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2057,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b00110010; c = 8'b10001101; // Expected: {'sum': 171, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b00110010; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2058,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00010110; c = 8'b11100110; // Expected: {'sum': 98, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00010110; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2059,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00001011; c = 8'b11011010; // Expected: {'sum': 113, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00001011; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2060,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00010101; c = 8'b10001100; // Expected: {'sum': 71, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00010101; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2061,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10011010; c = 8'b00000010; // Expected: {'sum': 13, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10011010; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2062,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b01101010; c = 8'b11101011; // Expected: {'sum': 230, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b01101010; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2063,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11010010; c = 8'b10001100; // Expected: {'sum': 0, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11010010; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2064,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11111100; c = 8'b10000110; // Expected: {'sum': 143, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11111100; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2065,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10011101; c = 8'b01101000; // Expected: {'sum': 9, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10011101; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2066,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b01011110; c = 8'b00110101; // Expected: {'sum': 67, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b01011110; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2067,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b10011100; c = 8'b11001010; // Expected: {'sum': 68, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b10011100; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2068,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11010101; c = 8'b00110001; // Expected: {'sum': 115, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11010101; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2069,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b10001010; c = 8'b10111110; // Expected: {'sum': 181, 'carry': 138}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b10001010; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2070,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b01100110; c = 8'b11000010; // Expected: {'sum': 108, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b01100110; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2071,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11111000; c = 8'b00100110; // Expected: {'sum': 189, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11111000; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2072,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11100111; c = 8'b11010101; // Expected: {'sum': 99, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11100111; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2073,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b11110101; c = 8'b00110000; // Expected: {'sum': 126, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b11110101; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2074,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11111110; c = 8'b11010001; // Expected: {'sum': 35, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11111110; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2075,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00100000; c = 8'b10001110; // Expected: {'sum': 169, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00100000; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2076,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b10000000; c = 8'b00100010; // Expected: {'sum': 8, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b10000000; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2077,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10111011; c = 8'b00011000; // Expected: {'sum': 197, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10111011; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2078,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10101000; c = 8'b11010111; // Expected: {'sum': 143, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10101000; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2079,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b10100100; c = 8'b00101010; // Expected: {'sum': 78, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b10100100; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2080,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b01110111; c = 8'b10111100; // Expected: {'sum': 126, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b01110111; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2081,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11010100; c = 8'b00110010; // Expected: {'sum': 195, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11010100; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2082,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b11000101; c = 8'b11100111; // Expected: {'sum': 121, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b11000101; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2083,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b01000110; c = 8'b00010001; // Expected: {'sum': 17, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b01000110; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2084,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00101111; c = 8'b01011101; // Expected: {'sum': 55, 'carry': 77}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00101111; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2085,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b00001000; c = 8'b11110110; // Expected: {'sum': 208, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b00001000; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2086,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b11001110; c = 8'b10000101; // Expected: {'sum': 144, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b11001110; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2087,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b11111100; c = 8'b11010010; // Expected: {'sum': 126, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b11111100; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2088,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b10000100; c = 8'b11101010; // Expected: {'sum': 243, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b10000100; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2089,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00100010; c = 8'b01011000; // Expected: {'sum': 143, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00100010; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2090,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b01100101; c = 8'b01100101; // Expected: {'sum': 182, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b01100101; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2091,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11010110; c = 8'b00111111; // Expected: {'sum': 205, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11010110; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2092,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11110111; c = 8'b00010101; // Expected: {'sum': 75, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11110111; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2093,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10000100; c = 8'b10011000; // Expected: {'sum': 132, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10000100; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2094,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b00111111; c = 8'b11001111; // Expected: {'sum': 96, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b00111111; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2095,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b00000100; c = 8'b00101100; // Expected: {'sum': 66, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b00000100; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2096,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b11100011; c = 8'b01111001; // Expected: {'sum': 174, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b11100011; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2097,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b00000010; c = 8'b11110111; // Expected: {'sum': 222, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b00000010; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2098,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10100100; c = 8'b11011000; // Expected: {'sum': 33, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10100100; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2099,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b00101000; c = 8'b10010011; // Expected: {'sum': 114, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b00101000; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b01100001; c = 8'b10101000; // Expected: {'sum': 167, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b01100001; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b01100010; c = 8'b10100011; // Expected: {'sum': 225, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b01100010; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b11111010; c = 8'b01011010; // Expected: {'sum': 159, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b11111010; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00001111; c = 8'b10001000; // Expected: {'sum': 58, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00001111; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00101111; c = 8'b01101000; // Expected: {'sum': 247, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00101111; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b00100100; c = 8'b11100111; // Expected: {'sum': 89, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b00100100; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b00111000; c = 8'b01101011; // Expected: {'sum': 182, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b00111000; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b00100001; c = 8'b11010111; // Expected: {'sum': 148, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b00100001; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00101001; c = 8'b00110010; // Expected: {'sum': 157, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00101001; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b11100011; c = 8'b11010010; // Expected: {'sum': 15, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b11100011; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11101000; c = 8'b11010001; // Expected: {'sum': 162, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11101000; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01101011; c = 8'b00101010; // Expected: {'sum': 148, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01101011; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00001110; c = 8'b11001101; // Expected: {'sum': 107, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00001110; c = 8'b11001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b00010010; c = 8'b10111000; // Expected: {'sum': 131, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b00010010; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b10100010; c = 8'b00010011; // Expected: {'sum': 78, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b10100010; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b10100101; c = 8'b01010000; // Expected: {'sum': 226, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b10100101; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b10010111; c = 8'b00010010; // Expected: {'sum': 117, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b10010111; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11011010; c = 8'b10010011; // Expected: {'sum': 158, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11011010; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10011110; c = 8'b11001101; // Expected: {'sum': 161, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10011110; c = 8'b11001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01101110; c = 8'b01001010; // Expected: {'sum': 47, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01101110; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11110010; c = 8'b11101110; // Expected: {'sum': 16, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11110010; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01010100; c = 8'b01110100; // Expected: {'sum': 163, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01010100; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01011100; c = 8'b00011100; // Expected: {'sum': 16, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01011100; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10010000; c = 8'b01111000; // Expected: {'sum': 146, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10010000; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b10111000; c = 8'b10001111; // Expected: {'sum': 90, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b10111000; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b10111100; c = 8'b11001111; // Expected: {'sum': 137, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b10111100; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01010000; c = 8'b10100101; // Expected: {'sum': 36, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01010000; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b11011101; c = 8'b10010011; // Expected: {'sum': 78, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b11011101; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11011010; c = 8'b10001111; // Expected: {'sum': 128, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11011010; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10100010; c = 8'b11001100; // Expected: {'sum': 11, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10100010; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b01001111; c = 8'b11110100; // Expected: {'sum': 198, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b01001111; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b01111101; c = 8'b11100000; // Expected: {'sum': 93, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b01111101; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11010001; c = 8'b00100100; // Expected: {'sum': 81, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11010001; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b11111001; c = 8'b00100100; // Expected: {'sum': 87, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b11111001; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b00000010; c = 8'b10111000; // Expected: {'sum': 86, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b00000010; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b00000101; c = 8'b01111111; // Expected: {'sum': 118, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b00000101; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b10001101; c = 8'b10100110; // Expected: {'sum': 251, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b10001101; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10100100; c = 8'b11001100; // Expected: {'sum': 85, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10100100; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b00110111; c = 8'b10011100; // Expected: {'sum': 180, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b00110111; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11111000; c = 8'b00100101; // Expected: {'sum': 138, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11111000; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b10101000; c = 8'b10010110; // Expected: {'sum': 61, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b10101000; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10111101; c = 8'b10111100; // Expected: {'sum': 250, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10111101; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00110011; c = 8'b01001010; // Expected: {'sum': 17, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00110011; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10000101; c = 8'b10011101; // Expected: {'sum': 104, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10000101; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b11000011; c = 8'b00101010; // Expected: {'sum': 174, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b11000011; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01000110; c = 8'b11001010; // Expected: {'sum': 139, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01000110; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10111110; c = 8'b01101100; // Expected: {'sum': 178, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10111110; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b00010000; c = 8'b10100110; // Expected: {'sum': 54, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b00010000; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00010010; c = 8'b11101011; // Expected: {'sum': 182, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00010010; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11010101; c = 8'b10101100; // Expected: {'sum': 106, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11010101; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 106, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00010100; c = 8'b01011010; // Expected: {'sum': 176, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00010100; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b00101100; c = 8'b01100110; // Expected: {'sum': 52, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b00101100; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10001101; c = 8'b01110000; // Expected: {'sum': 105, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10001101; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10011001; c = 8'b00001110; // Expected: {'sum': 155, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10011001; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10110101; c = 8'b11110110; // Expected: {'sum': 221, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10110101; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01001110; c = 8'b00010011; // Expected: {'sum': 193, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01001110; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b01001101; c = 8'b11001001; // Expected: {'sum': 10, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b01001101; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00100011; c = 8'b00001101; // Expected: {'sum': 37, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00100011; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10010110; c = 8'b11111001; // Expected: {'sum': 254, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10010110; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b01010111; c = 8'b00000010; // Expected: {'sum': 118, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b01010111; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b11101001; c = 8'b00000100; // Expected: {'sum': 198, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b11101001; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01111000; c = 8'b01011011; // Expected: {'sum': 191, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01111000; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b10111001; c = 8'b00111000; // Expected: {'sum': 14, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b10111001; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10111101; c = 8'b10100111; // Expected: {'sum': 0, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10111101; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b10000010; c = 8'b01001010; // Expected: {'sum': 77, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b10000010; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b11101000; c = 8'b10011001; // Expected: {'sum': 91, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b11101000; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00000100; c = 8'b00111011; // Expected: {'sum': 180, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00000100; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00111000; c = 8'b10000011; // Expected: {'sum': 20, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00111000; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00110011; c = 8'b00111110; // Expected: {'sum': 147, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00110011; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10011000; c = 8'b10010011; // Expected: {'sum': 113, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10011000; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11101100; c = 8'b10000101; // Expected: {'sum': 213, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11101100; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b10010100; c = 8'b11000000; // Expected: {'sum': 140, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b10010100; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01011001; c = 8'b01001001; // Expected: {'sum': 147, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01011001; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01101001; c = 8'b01111010; // Expected: {'sum': 143, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01101001; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10000001; c = 8'b11111100; // Expected: {'sum': 177, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10000001; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b11101110; c = 8'b00111100; // Expected: {'sum': 181, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b11101110; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b11011101; c = 8'b01001011; // Expected: {'sum': 203, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b11011101; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b10011101; c = 8'b10001001; // Expected: {'sum': 6, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b10011101; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b00010010; c = 8'b11001110; // Expected: {'sum': 24, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b00010010; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00111000; c = 8'b10111101; // Expected: {'sum': 143, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00111000; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10010000; c = 8'b01011110; // Expected: {'sum': 182, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10010000; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b11100100; c = 8'b01101011; // Expected: {'sum': 66, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b11100100; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01111011; c = 8'b11011110; // Expected: {'sum': 159, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01111011; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00010100; c = 8'b11100101; // Expected: {'sum': 130, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00010100; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01010011; c = 8'b11000001; // Expected: {'sum': 52, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01010011; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b01010101; c = 8'b10011000; // Expected: {'sum': 185, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b01010101; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10011101; c = 8'b01010011; // Expected: {'sum': 162, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10011101; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10001100; c = 8'b01011110; // Expected: {'sum': 195, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10001100; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b00011100; c = 8'b11011110; // Expected: {'sum': 27, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b00011100; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11011011; c = 8'b10000110; // Expected: {'sum': 94, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11011011; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b11010110; c = 8'b00100000; // Expected: {'sum': 147, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b11010110; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10100000; c = 8'b11011100; // Expected: {'sum': 136, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10100000; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01111111; c = 8'b10010000; // Expected: {'sum': 177, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01111111; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11000101; c = 8'b00100010; // Expected: {'sum': 53, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11000101; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00001110; c = 8'b10110000; // Expected: {'sum': 44, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00001110; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b10110111; c = 8'b10111111; // Expected: {'sum': 164, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b10110111; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b00001011; c = 8'b11101010; // Expected: {'sum': 248, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b00001011; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01011110; c = 8'b11110111; // Expected: {'sum': 202, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01011110; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b00010011; c = 8'b10001110; // Expected: {'sum': 63, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b00010011; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01110010; c = 8'b10010101; // Expected: {'sum': 139, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01110010; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11110100; c = 8'b10000111; // Expected: {'sum': 250, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11110100; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11100100; c = 8'b10111110; // Expected: {'sum': 191, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11100100; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10011110; c = 8'b01010001; // Expected: {'sum': 157, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10011110; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00001100; c = 8'b11011110; // Expected: {'sum': 159, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00001100; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01111000; c = 8'b10110010; // Expected: {'sum': 22, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01111000; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10101110; c = 8'b01110000; // Expected: {'sum': 58, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10101110; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10010100; c = 8'b00000100; // Expected: {'sum': 84, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10010100; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10110100; c = 8'b10100100; // Expected: {'sum': 48, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10110100; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00011111; c = 8'b01011111; // Expected: {'sum': 7, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00011111; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11110110; c = 8'b10000100; // Expected: {'sum': 217, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11110110; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01101110; c = 8'b01101100; // Expected: {'sum': 95, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01101110; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b01101101; c = 8'b11011001; // Expected: {'sum': 230, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b01101101; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00000110; c = 8'b10010111; // Expected: {'sum': 27, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00000110; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00010010; c = 8'b00001011; // Expected: {'sum': 112, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00010010; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11001100; c = 8'b01111110; // Expected: {'sum': 142, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11001100; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b11100111; c = 8'b00010000; // Expected: {'sum': 140, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b11100111; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b00110011; c = 8'b01111101; // Expected: {'sum': 6, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b00110011; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b00100001; c = 8'b00101011; // Expected: {'sum': 157, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b00100001; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b01000111; c = 8'b11011110; // Expected: {'sum': 215, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b01000111; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01011001; c = 8'b11100101; // Expected: {'sum': 105, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01011001; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10010001; c = 8'b10110000; // Expected: {'sum': 186, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10010001; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10100011; c = 8'b10101101; // Expected: {'sum': 32, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10100011; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b01101110; c = 8'b11111101; // Expected: {'sum': 22, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b01101110; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b00100001; c = 8'b10100110; // Expected: {'sum': 74, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b00100001; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b10000100; c = 8'b00000111; // Expected: {'sum': 19, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b10000100; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b00010111; c = 8'b11110011; // Expected: {'sum': 18, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b00010111; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01100001; c = 8'b01011100; // Expected: {'sum': 216, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01100001; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10011111; c = 8'b11101100; // Expected: {'sum': 54, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10011111; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00011001; c = 8'b01000011; // Expected: {'sum': 144, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00011001; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01111100; c = 8'b01111111; // Expected: {'sum': 138, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01111100; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b10101111; c = 8'b00110001; // Expected: {'sum': 254, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b10101111; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b11000110; c = 8'b00110110; // Expected: {'sum': 192, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b11000110; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b00001101; c = 8'b00000111; // Expected: {'sum': 90, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b00001101; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b01110010; c = 8'b01010110; // Expected: {'sum': 213, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b01110010; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11011000; c = 8'b00010110; // Expected: {'sum': 75, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11011000; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01100101; c = 8'b10110100; // Expected: {'sum': 214, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01100101; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11001101; c = 8'b11110101; // Expected: {'sum': 115, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11001101; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10001011; c = 8'b01110101; // Expected: {'sum': 252, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10001011; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10011001; c = 8'b10011100; // Expected: {'sum': 65, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10011001; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01010110; c = 8'b01010010; // Expected: {'sum': 156, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01010110; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11101110; c = 8'b01001010; // Expected: {'sum': 178, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11101110; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00001011; c = 8'b00101011; // Expected: {'sum': 72, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00001011; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b11000011; c = 8'b01100100; // Expected: {'sum': 215, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b11000011; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00010101; c = 8'b01010101; // Expected: {'sum': 65, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00010101; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11000001; c = 8'b01110110; // Expected: {'sum': 103, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11000001; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11010011; c = 8'b11011111; // Expected: {'sum': 137, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11010011; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11110011; c = 8'b10111000; // Expected: {'sum': 39, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11110011; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10001110; c = 8'b00110011; // Expected: {'sum': 172, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10001110; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00010100; c = 8'b11101111; // Expected: {'sum': 160, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00010100; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11110111; c = 8'b01011100; // Expected: {'sum': 95, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11110111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11011101; c = 8'b00011001; // Expected: {'sum': 6, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11011101; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10001110; c = 8'b01111000; // Expected: {'sum': 215, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10001110; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b01101011; c = 8'b11001011; // Expected: {'sum': 252, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b01101011; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11000011; c = 8'b11011001; // Expected: {'sum': 216, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11000011; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00100001; c = 8'b01000111; // Expected: {'sum': 154, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00100001; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00101100; c = 8'b00010100; // Expected: {'sum': 116, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00101100; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b11011010; c = 8'b01001101; // Expected: {'sum': 213, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b11011010; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11110101; c = 8'b10101111; // Expected: {'sum': 130, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11110101; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00011111; c = 8'b10001111; // Expected: {'sum': 63, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00011111; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00001101; c = 8'b00100101; // Expected: {'sum': 150, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00001101; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b11000011; c = 8'b01110000; // Expected: {'sum': 120, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b11000011; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10011010; c = 8'b00111001; // Expected: {'sum': 187, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10011010; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00111001; c = 8'b11010001; // Expected: {'sum': 206, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00111001; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10010111; c = 8'b00001010; // Expected: {'sum': 248, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10010111; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b00000011; c = 8'b00110000; // Expected: {'sum': 242, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b00000011; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01100111; c = 8'b01011100; // Expected: {'sum': 210, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01100111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b00110100; c = 8'b10110111; // Expected: {'sum': 148, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b00110100; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10000111; c = 8'b00010101; // Expected: {'sum': 96, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10000111; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b10111000; c = 8'b00111101; // Expected: {'sum': 132, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b10111000; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10100111; c = 8'b11110101; // Expected: {'sum': 202, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10100111; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00010011; c = 8'b10111000; // Expected: {'sum': 48, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00010011; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b10111110; c = 8'b00010011; // Expected: {'sum': 24, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b10111110; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 24, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10100101; c = 8'b11100111; // Expected: {'sum': 8, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10100101; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b00101001; c = 8'b10100110; // Expected: {'sum': 191, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b00101001; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10101010; c = 8'b01100001; // Expected: {'sum': 20, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10101010; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01100000; c = 8'b01111001; // Expected: {'sum': 159, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01100000; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01011001; c = 8'b01110100; // Expected: {'sum': 148, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01011001; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b11110100; c = 8'b11010101; // Expected: {'sum': 21, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b11110100; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01000100; c = 8'b00111010; // Expected: {'sum': 253, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01000100; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b10100010; c = 8'b10011001; // Expected: {'sum': 25, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b10100010; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11010000; c = 8'b01000110; // Expected: {'sum': 246, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11010000; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10100101; c = 8'b11001000; // Expected: {'sum': 32, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10100101; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10110111; c = 8'b01111111; // Expected: {'sum': 11, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10110111; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b11010001; c = 8'b00001110; // Expected: {'sum': 53, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b11010001; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b00001010; c = 8'b01001111; // Expected: {'sum': 25, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b00001010; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00111101; c = 8'b01000100; // Expected: {'sum': 135, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00111101; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10010011; c = 8'b11001011; // Expected: {'sum': 226, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10010011; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10101100; c = 8'b10101011; // Expected: {'sum': 101, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10101100; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b10011011; c = 8'b00110010; // Expected: {'sum': 127, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b10011011; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00101011; c = 8'b01100000; // Expected: {'sum': 54, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00101011; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01000001; c = 8'b11011111; // Expected: {'sum': 145, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01000001; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b10001001; c = 8'b01000010; // Expected: {'sum': 145, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b10001001; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10100010; c = 8'b11011001; // Expected: {'sum': 188, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10100010; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b01101010; c = 8'b01011000; // Expected: {'sum': 46, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b01101010; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11001111; c = 8'b00101010; // Expected: {'sum': 37, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11001111; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b11000011; c = 8'b11101000; // Expected: {'sum': 135, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b11000011; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b11000000; c = 8'b11001111; // Expected: {'sum': 215, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b11000000; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b01110100; c = 8'b00000110; // Expected: {'sum': 219, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b01110100; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b11000101; c = 8'b11111110; // Expected: {'sum': 246, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b11000101; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b00110100; c = 8'b00011111; // Expected: {'sum': 78, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b00110100; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b00000110; c = 8'b11100000; // Expected: {'sum': 38, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b00000110; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b01011100; c = 8'b01001000; // Expected: {'sum': 186, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b01011100; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10011010; c = 8'b00100011; // Expected: {'sum': 245, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10011010; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b00000001; c = 8'b10111100; // Expected: {'sum': 123, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b00000001; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10001100; c = 8'b10011100; // Expected: {'sum': 236, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10001100; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b11110111; c = 8'b00011010; // Expected: {'sum': 163, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b11110111; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00101110; c = 8'b01111101; // Expected: {'sum': 197, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00101110; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b11100101; c = 8'b11100110; // Expected: {'sum': 144, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b11100101; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b11110101; c = 8'b00111101; // Expected: {'sum': 34, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b11110101; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10100010; c = 8'b00001100; // Expected: {'sum': 229, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10100010; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b00001101; c = 8'b00011010; // Expected: {'sum': 94, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b00001101; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b10011010; c = 8'b00110110; // Expected: {'sum': 255, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b10011010; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10011100; c = 8'b01010001; // Expected: {'sum': 241, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10011100; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b10111111; c = 8'b01011010; // Expected: {'sum': 29, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b10111111; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01101110; c = 8'b00010011; // Expected: {'sum': 55, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01101110; c = 8'b00010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00010001; c = 8'b11000111; // Expected: {'sum': 141, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00010001; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b00010100; c = 8'b10101000; // Expected: {'sum': 143, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b00010100; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b11001011; c = 8'b01111001; // Expected: {'sum': 45, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b11001011; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01101100; c = 8'b01010011; // Expected: {'sum': 154, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01101100; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10111100; c = 8'b00001000; // Expected: {'sum': 136, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10111100; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00101001; c = 8'b00101111; // Expected: {'sum': 55, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00101001; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00011110; c = 8'b00001100; // Expected: {'sum': 95, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00011110; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b01100010; c = 8'b10111110; // Expected: {'sum': 89, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b01100010; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b00011100; c = 8'b00011011; // Expected: {'sum': 100, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b00011100; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01111111; c = 8'b11010010; // Expected: {'sum': 124, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01111111; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10100110; c = 8'b11001111; // Expected: {'sum': 50, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10100110; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10101100; c = 8'b00100110; // Expected: {'sum': 240, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10101100; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00010000; c = 8'b10001010; // Expected: {'sum': 251, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00010000; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b10001011; c = 8'b11001001; // Expected: {'sum': 76, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b10001011; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01011000; c = 8'b10100100; // Expected: {'sum': 147, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01011000; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11101001; c = 8'b11001100; // Expected: {'sum': 209, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11101001; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b01101011; c = 8'b01101001; // Expected: {'sum': 232, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b01101011; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00111011; c = 8'b01101010; // Expected: {'sum': 77, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00111011; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11100100; c = 8'b10101101; // Expected: {'sum': 192, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11100100; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11100110; c = 8'b11100110; // Expected: {'sum': 22, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11100110; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11100011; c = 8'b10001110; // Expected: {'sum': 223, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11100011; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b00101110; c = 8'b01011101; // Expected: {'sum': 235, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b00101110; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b01000111; c = 8'b01110001; // Expected: {'sum': 102, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b01000111; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10100110; c = 8'b10010011; // Expected: {'sum': 15, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10100110; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01000001; c = 8'b10000001; // Expected: {'sum': 179, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01000001; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10100001; c = 8'b10011010; // Expected: {'sum': 103, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10100001; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10100101; c = 8'b00111010; // Expected: {'sum': 67, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10100101; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01001001; c = 8'b01101110; // Expected: {'sum': 38, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01001001; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b11000111; c = 8'b10111001; // Expected: {'sum': 162, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b11000111; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11101000; c = 8'b10011110; // Expected: {'sum': 206, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11101000; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11100000; c = 8'b00000000; // Expected: {'sum': 63, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11100000; c = 8'b00000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01100110; c = 8'b10010000; // Expected: {'sum': 89, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01100110; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10011101; c = 8'b10011010; // Expected: {'sum': 191, 'carry': 152}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10011101; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01001100; c = 8'b00110000; // Expected: {'sum': 241, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01001100; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b11100010; c = 8'b00100010; // Expected: {'sum': 205, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b11100010; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11000000; c = 8'b00001011; // Expected: {'sum': 62, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11000000; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b11110010; c = 8'b00111100; // Expected: {'sum': 111, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b11110010; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10011110; c = 8'b01000111; // Expected: {'sum': 143, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10011110; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b11100110; c = 8'b10101001; // Expected: {'sum': 104, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b11100110; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b10001110; c = 8'b11110101; // Expected: {'sum': 26, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b10001110; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01000001; c = 8'b10110111; // Expected: {'sum': 105, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01000001; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10111010; c = 8'b11011011; // Expected: {'sum': 250, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10111010; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b11011111; c = 8'b11000100; // Expected: {'sum': 199, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b11011111; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10100011; c = 8'b01010110; // Expected: {'sum': 92, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10100011; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10101010; c = 8'b01100110; // Expected: {'sum': 174, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10101010; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00111100; c = 8'b11001001; // Expected: {'sum': 27, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00111100; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 27, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01001100; c = 8'b10101000; // Expected: {'sum': 85, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01001100; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10000110; c = 8'b10110100; // Expected: {'sum': 43, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10000110; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b10101001; c = 8'b01101011; // Expected: {'sum': 138, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b10101001; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00010001; c = 8'b10010100; // Expected: {'sum': 143, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00010001; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b11100010; c = 8'b01001000; // Expected: {'sum': 101, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b11100010; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b11110011; c = 8'b00000001; // Expected: {'sum': 113, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b11110011; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01101001; c = 8'b00011111; // Expected: {'sum': 254, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01101001; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b11110001; c = 8'b00010101; // Expected: {'sum': 43, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b11110001; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11001110; c = 8'b10010011; // Expected: {'sum': 35, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11001110; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01010000; c = 8'b00011101; // Expected: {'sum': 169, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01010000; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11011000; c = 8'b01011100; // Expected: {'sum': 166, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11011000; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b00101100; c = 8'b11110100; // Expected: {'sum': 135, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b00101100; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b00000011; c = 8'b00100100; // Expected: {'sum': 87, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b00000011; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b01100000; c = 8'b11011000; // Expected: {'sum': 169, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b01100000; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b11111011; c = 8'b10101110; // Expected: {'sum': 76, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b11111011; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b10000000; c = 8'b00100011; // Expected: {'sum': 159, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b10000000; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00110101; c = 8'b11101111; // Expected: {'sum': 169, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00110101; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01110000; c = 8'b01010100; // Expected: {'sum': 44, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01110000; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11100110; c = 8'b11011010; // Expected: {'sum': 75, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11100110; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b11101111; c = 8'b00110011; // Expected: {'sum': 110, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b11101111; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11011101; c = 8'b10001100; // Expected: {'sum': 250, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11011101; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11011000; c = 8'b00110010; // Expected: {'sum': 10, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11011000; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00011000; c = 8'b10101101; // Expected: {'sum': 132, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00011000; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11100110; c = 8'b00001010; // Expected: {'sum': 155, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11100110; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10010110; c = 8'b00110001; // Expected: {'sum': 241, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10010110; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10001000; c = 8'b01011100; // Expected: {'sum': 107, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10001000; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b00010011; c = 8'b01110000; // Expected: {'sum': 98, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b00010011; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00101010; c = 8'b10000001; // Expected: {'sum': 233, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00101010; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11010101; c = 8'b01010000; // Expected: {'sum': 155, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11010101; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b01011011; c = 8'b01010010; // Expected: {'sum': 245, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b01011011; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b01011110; c = 8'b11001101; // Expected: {'sum': 45, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b01011110; c = 8'b11001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10101101; c = 8'b01011110; // Expected: {'sum': 191, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10101101; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00010000; c = 8'b10100010; // Expected: {'sum': 158, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00010000; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b11111110; c = 8'b11011100; // Expected: {'sum': 216, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b11111110; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01001111; c = 8'b10110001; // Expected: {'sum': 11, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01001111; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01101111; c = 8'b00000110; // Expected: {'sum': 109, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01101111; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b11110110; c = 8'b10000011; // Expected: {'sum': 240, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b11110110; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10001000; c = 8'b01110110; // Expected: {'sum': 198, 'carry': 56}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10001000; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01010001; c = 8'b10100001; // Expected: {'sum': 55, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01010001; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10100011; c = 8'b00100111; // Expected: {'sum': 153, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10100011; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b11101101; c = 8'b10110100; // Expected: {'sum': 109, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b11101101; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10000011; c = 8'b00010000; // Expected: {'sum': 41, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10000011; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11101000; c = 8'b01101101; // Expected: {'sum': 208, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11101000; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10011011; c = 8'b01000001; // Expected: {'sum': 255, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10011011; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11110101; c = 8'b01011100; // Expected: {'sum': 93, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11110101; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b00001011; c = 8'b10101100; // Expected: {'sum': 223, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b00001011; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b11011011; c = 8'b11111001; // Expected: {'sum': 130, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b11011011; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10111111; c = 8'b00111011; // Expected: {'sum': 186, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10111111; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b11000111; c = 8'b00110000; // Expected: {'sum': 31, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b11000111; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b11101100; c = 8'b00100101; // Expected: {'sum': 73, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b11101100; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b10000111; c = 8'b10000101; // Expected: {'sum': 22, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b10000111; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10101110; c = 8'b10100110; // Expected: {'sum': 16, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10101110; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01110000; c = 8'b10000011; // Expected: {'sum': 238, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01110000; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01010111; c = 8'b10100100; // Expected: {'sum': 58, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01010111; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01111001; c = 8'b11100100; // Expected: {'sum': 194, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01111001; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b00111100; c = 8'b01110001; // Expected: {'sum': 116, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b00111100; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b01011110; c = 8'b10011101; // Expected: {'sum': 140, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b01011110; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11000111; c = 8'b01011101; // Expected: {'sum': 30, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11000111; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b10101111; c = 8'b11111011; // Expected: {'sum': 215, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b10101111; c = 8'b11111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b11100101; c = 8'b10110101; // Expected: {'sum': 202, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b11100101; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b11100010; c = 8'b01000101; // Expected: {'sum': 165, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b11100010; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01111011; c = 8'b10010000; // Expected: {'sum': 20, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01111011; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11101001; c = 8'b10011100; // Expected: {'sum': 8, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11101001; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b00111110; c = 8'b00010010; // Expected: {'sum': 120, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b00111110; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10011000; c = 8'b00101101; // Expected: {'sum': 21, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10011000; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10100001; c = 8'b11110001; // Expected: {'sum': 182, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10100001; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b00001110; c = 8'b10100111; // Expected: {'sum': 49, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b00001110; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b10101011; c = 8'b00101111; // Expected: {'sum': 44, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b10101011; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01011110; c = 8'b11010110; // Expected: {'sum': 143, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01011110; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10011101; c = 8'b01001001; // Expected: {'sum': 32, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10011101; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b11100000; c = 8'b11000010; // Expected: {'sum': 32, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b11100000; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b10111011; c = 8'b01100111; // Expected: {'sum': 73, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b10111011; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b00101000; c = 8'b01011100; // Expected: {'sum': 110, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b00101000; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b10110110; c = 8'b11110001; // Expected: {'sum': 173, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b10110110; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11101001; c = 8'b00110000; // Expected: {'sum': 37, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11101001; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01001011; c = 8'b00010101; // Expected: {'sum': 1, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01001011; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10010001; c = 8'b10101010; // Expected: {'sum': 252, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10010001; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 252, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10111011; c = 8'b01101000; // Expected: {'sum': 232, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10111011; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b00010100; c = 8'b11000100; // Expected: {'sum': 108, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b00010100; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b11000000; c = 8'b01001111; // Expected: {'sum': 113, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b11000000; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b00101110; c = 8'b10100010; // Expected: {'sum': 174, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b00101110; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00010111; c = 8'b01010100; // Expected: {'sum': 101, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00010111; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01101000; c = 8'b01101110; // Expected: {'sum': 195, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01101000; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b00100111; c = 8'b10111011; // Expected: {'sum': 9, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b00100111; c = 8'b10111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b10111101; c = 8'b00101101; // Expected: {'sum': 186, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b10111101; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01001100; c = 8'b10110010; // Expected: {'sum': 212, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01001100; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b10100101; c = 8'b01001001; // Expected: {'sum': 138, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b10100101; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01001110; c = 8'b10101101; // Expected: {'sum': 156, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01001110; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b10111000; c = 8'b00100001; // Expected: {'sum': 69, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b10111000; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00110110; c = 8'b01101100; // Expected: {'sum': 234, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00110110; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11001100; c = 8'b00111000; // Expected: {'sum': 158, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11001100; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b11111100; c = 8'b01010010; // Expected: {'sum': 123, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b11111100; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b10101010; c = 8'b01000001; // Expected: {'sum': 49, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b10101010; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b00001001; c = 8'b10010101; // Expected: {'sum': 78, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b00001001; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b11100001; c = 8'b10001101; // Expected: {'sum': 147, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b11100001; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b00010001; c = 8'b00111000; // Expected: {'sum': 68, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b00010001; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b11110100; c = 8'b00110011; // Expected: {'sum': 72, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b11110100; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b11011001; c = 8'b10010110; // Expected: {'sum': 134, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b11011001; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11101101; c = 8'b01010100; // Expected: {'sum': 43, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11101101; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b01100110; c = 8'b11101010; // Expected: {'sum': 200, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b01100110; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10101100; c = 8'b00110110; // Expected: {'sum': 11, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10101100; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b10101111; c = 8'b01111011; // Expected: {'sum': 223, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b10101111; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10000010; c = 8'b00111000; // Expected: {'sum': 253, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10000010; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10111110; c = 8'b00101010; // Expected: {'sum': 146, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10111110; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b00101011; c = 8'b10101011; // Expected: {'sum': 191, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b00101011; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b11101011; c = 8'b11010011; // Expected: {'sum': 181, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b11101011; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10000111; c = 8'b01001011; // Expected: {'sum': 103, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10000111; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10111101; c = 8'b11001111; // Expected: {'sum': 137, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10111101; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00011010; c = 8'b10010011; // Expected: {'sum': 131, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00011010; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b11011001; c = 8'b01111001; // Expected: {'sum': 216, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b11011001; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10011101; c = 8'b11111010; // Expected: {'sum': 131, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10011101; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10101101; c = 8'b01010110; // Expected: {'sum': 165, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10101101; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b11001101; c = 8'b10110110; // Expected: {'sum': 73, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b11001101; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00110001; c = 8'b00000010; // Expected: {'sum': 237, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00110001; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b01100010; c = 8'b10000111; // Expected: {'sum': 109, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b01100010; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11111010; c = 8'b01111001; // Expected: {'sum': 185, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11111010; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b01011001; c = 8'b00001101; // Expected: {'sum': 164, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b01011001; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b11101000; c = 8'b01001001; // Expected: {'sum': 113, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b11101000; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00100010; c = 8'b01100010; // Expected: {'sum': 51, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00100010; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01110010; c = 8'b11010011; // Expected: {'sum': 79, 'carry': 242}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01110010; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01111111; c = 8'b00011100; // Expected: {'sum': 245, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01111111; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b00001100; c = 8'b01000001; // Expected: {'sum': 51, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b00001100; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11101110; c = 8'b00001010; // Expected: {'sum': 236, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11101110; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00010011; c = 8'b11011001; // Expected: {'sum': 133, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00010011; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 133, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00100011; c = 8'b11001011; // Expected: {'sum': 83, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00100011; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10110100; c = 8'b01111101; // Expected: {'sum': 41, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10110100; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b01100100; c = 8'b01011110; // Expected: {'sum': 6, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b01100100; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10111100; c = 8'b11111001; // Expected: {'sum': 104, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10111100; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b10010001; c = 8'b00000111; // Expected: {'sum': 205, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b10010001; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00110001; c = 8'b00110010; // Expected: {'sum': 50, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00110001; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10101001; c = 8'b01111100; // Expected: {'sum': 218, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10101001; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b00110011; c = 8'b01001010; // Expected: {'sum': 145, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b00110011; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b10111000; c = 8'b01111111; // Expected: {'sum': 189, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b10111000; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b01100110; c = 8'b11000101; // Expected: {'sum': 198, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b01100110; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b10111110; c = 8'b00100000; // Expected: {'sum': 123, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b10111110; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10000000; c = 8'b10110110; // Expected: {'sum': 94, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10000000; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00011101; c = 8'b01111000; // Expected: {'sum': 149, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00011101; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01111010; c = 8'b11011101; // Expected: {'sum': 48, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01111010; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11100100; c = 8'b01010000; // Expected: {'sum': 165, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11100100; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01100011; c = 8'b01000110; // Expected: {'sum': 12, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01100011; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01101011; c = 8'b01011000; // Expected: {'sum': 163, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01101011; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00010110; c = 8'b00001011; // Expected: {'sum': 70, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00010110; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00001111; c = 8'b01001101; // Expected: {'sum': 226, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00001111; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b00011001; c = 8'b10101001; // Expected: {'sum': 154, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b00011001; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00101111; c = 8'b11011011; // Expected: {'sum': 244, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00101111; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11011000; c = 8'b00000101; // Expected: {'sum': 244, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11011000; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 244, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b10110011; c = 8'b00011111; // Expected: {'sum': 172, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b10110011; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11010110; c = 8'b10010110; // Expected: {'sum': 115, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11010110; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 115, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b01010001; c = 8'b01100100; // Expected: {'sum': 49, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b01010001; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b10100110; c = 8'b10101001; // Expected: {'sum': 112, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b10100110; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01010111; c = 8'b11110101; // Expected: {'sum': 143, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01010111; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b10100011; c = 8'b10001110; // Expected: {'sum': 79, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b10100011; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01111001; c = 8'b01000111; // Expected: {'sum': 205, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01111001; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11100010; c = 8'b10100001; // Expected: {'sum': 144, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11100010; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00110100; c = 8'b10011100; // Expected: {'sum': 160, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00110100; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b01111011; c = 8'b10000011; // Expected: {'sum': 48, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b01111011; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b11001011; c = 8'b00101101; // Expected: {'sum': 5, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b11001011; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01010101; c = 8'b00110000; // Expected: {'sum': 212, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01010101; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10000111; c = 8'b11110000; // Expected: {'sum': 127, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10000111; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01101101; c = 8'b01010110; // Expected: {'sum': 254, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01101101; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10101011; c = 8'b10011111; // Expected: {'sum': 240, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10101011; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b00000001; c = 8'b01101111; // Expected: {'sum': 141, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b00000001; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10011010; c = 8'b10111111; // Expected: {'sum': 196, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10011010; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b10111110; c = 8'b01000000; // Expected: {'sum': 236, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b10111110; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b10110100; c = 8'b10110010; // Expected: {'sum': 134, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b10110100; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00001110; c = 8'b10101011; // Expected: {'sum': 95, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00001110; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10101000; c = 8'b11100001; // Expected: {'sum': 64, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10101000; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01100110; c = 8'b00100101; // Expected: {'sum': 206, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01100110; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10100011; c = 8'b01111000; // Expected: {'sum': 82, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10100011; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b01011001; c = 8'b00010101; // Expected: {'sum': 211, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b01011001; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10000100; c = 8'b10011100; // Expected: {'sum': 188, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10000100; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10011100; c = 8'b11100110; // Expected: {'sum': 142, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10011100; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00011110; c = 8'b01100001; // Expected: {'sum': 128, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00011110; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b00011001; c = 8'b11010011; // Expected: {'sum': 238, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b00011001; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b11110110; c = 8'b10110110; // Expected: {'sum': 180, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b11110110; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b00111100; c = 8'b00111100; // Expected: {'sum': 233, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b00111100; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00001010; c = 8'b00001110; // Expected: {'sum': 125, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00001010; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01000101; c = 8'b01110101; // Expected: {'sum': 159, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01000101; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b00011100; c = 8'b11100010; // Expected: {'sum': 145, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b00011100; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b01100011; c = 8'b10101110; // Expected: {'sum': 86, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b01100011; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b10000000; c = 8'b11110100; // Expected: {'sum': 106, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b10000000; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 106, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b11111100; c = 8'b11101110; // Expected: {'sum': 233, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b11111100; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00000111; c = 8'b10101111; // Expected: {'sum': 41, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00000111; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11000110; c = 8'b00001110; // Expected: {'sum': 89, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11000110; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b00101001; c = 8'b10001110; // Expected: {'sum': 19, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b00101001; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10110011; c = 8'b00000110; // Expected: {'sum': 8, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10110011; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10001110; c = 8'b01011001; // Expected: {'sum': 154, 'carry': 77}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10001110; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b10111010; c = 8'b01001110; // Expected: {'sum': 98, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b10111010; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01111111; c = 8'b11010001; // Expected: {'sum': 202, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01111111; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b00011000; c = 8'b01001000; // Expected: {'sum': 107, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b00011000; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01011110; c = 8'b01001100; // Expected: {'sum': 246, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01011110; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01101001; c = 8'b10100010; // Expected: {'sum': 123, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01101001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b01010000; c = 8'b11010101; // Expected: {'sum': 0, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b01010000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11110101; c = 8'b01111000; // Expected: {'sum': 108, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11110101; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b10111100; c = 8'b11010010; // Expected: {'sum': 216, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b10111100; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b10010011; c = 8'b01101101; // Expected: {'sum': 191, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b10010011; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b10111101; c = 8'b00101111; // Expected: {'sum': 41, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b10111101; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01110010; c = 8'b00101011; // Expected: {'sum': 241, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01110010; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01101110; c = 8'b01011000; // Expected: {'sum': 74, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01101110; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b01111011; c = 8'b01101100; // Expected: {'sum': 40, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b01111011; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b00111011; c = 8'b01111101; // Expected: {'sum': 43, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b00111011; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b10101111; c = 8'b00110100; // Expected: {'sum': 239, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b10101111; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b10001010; c = 8'b11101011; // Expected: {'sum': 5, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b10001010; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00101000; c = 8'b11011000; // Expected: {'sum': 180, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00101000; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b00011110; c = 8'b01001000; // Expected: {'sum': 2, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b00011110; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01010010; c = 8'b11000010; // Expected: {'sum': 160, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01010010; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b01101010; c = 8'b01110000; // Expected: {'sum': 63, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b01101010; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b10001111; c = 8'b01100001; // Expected: {'sum': 195, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b10001111; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b10110000; c = 8'b10111001; // Expected: {'sum': 22, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b10110000; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10011000; c = 8'b11100101; // Expected: {'sum': 181, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10011000; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11101110; c = 8'b01000001; // Expected: {'sum': 50, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11101110; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01101010; c = 8'b01110000; // Expected: {'sum': 121, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01101010; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10101101; c = 8'b10010101; // Expected: {'sum': 50, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10101101; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b00000000; c = 8'b00000110; // Expected: {'sum': 88, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b00000000; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00111111; c = 8'b00100000; // Expected: {'sum': 129, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00111111; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11101100; c = 8'b10010111; // Expected: {'sum': 216, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11101100; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b01000111; c = 8'b11000100; // Expected: {'sum': 153, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b01000111; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b00101110; c = 8'b00011101; // Expected: {'sum': 121, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b00101110; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b11011110; c = 8'b00000110; // Expected: {'sum': 211, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b11011110; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01000010; c = 8'b11100011; // Expected: {'sum': 74, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01000010; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b11011000; c = 8'b01011100; // Expected: {'sum': 114, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b11011000; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11010110; c = 8'b10010000; // Expected: {'sum': 19, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11010110; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b01100100; c = 8'b01010001; // Expected: {'sum': 14, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b01100100; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b11011010; c = 8'b11111111; // Expected: {'sum': 32, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b11011010; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10100000; c = 8'b11110000; // Expected: {'sum': 95, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10100000; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b00111100; c = 8'b11100101; // Expected: {'sum': 155, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b00111100; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11001100; c = 8'b01100000; // Expected: {'sum': 93, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11001100; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10001101; c = 8'b00101100; // Expected: {'sum': 187, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10001101; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01110101; c = 8'b10110111; // Expected: {'sum': 169, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01110101; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11110101; c = 8'b00110111; // Expected: {'sum': 107, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11110101; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10101111; c = 8'b10110010; // Expected: {'sum': 169, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10101111; c = 8'b10110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10111001; c = 8'b11110111; // Expected: {'sum': 161, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10111001; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b11110110; c = 8'b11000100; // Expected: {'sum': 74, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b11110110; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11110001; c = 8'b10001111; // Expected: {'sum': 143, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11110001; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b01001001; c = 8'b00001001; // Expected: {'sum': 36, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b01001001; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b11111001; c = 8'b10111001; // Expected: {'sum': 165, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b11111001; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b00110110; c = 8'b01100110; // Expected: {'sum': 218, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b00110110; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b10101001; c = 8'b01011010; // Expected: {'sum': 81, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b10101001; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b00110000; c = 8'b01001001; // Expected: {'sum': 178, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b00110000; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b11101011; c = 8'b11101001; // Expected: {'sum': 140, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b11101011; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b01101110; c = 8'b10111001; // Expected: {'sum': 91, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b01101110; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10100111; c = 8'b00100100; // Expected: {'sum': 223, 'carry': 36}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10100111; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b00101100; c = 8'b11001111; // Expected: {'sum': 98, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b00101100; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11101101; c = 8'b01000111; // Expected: {'sum': 160, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11101101; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00111110; c = 8'b10011001; // Expected: {'sum': 10, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00111110; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b00100000; c = 8'b01100111; // Expected: {'sum': 14, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b00100000; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b00100000; c = 8'b11110110; // Expected: {'sum': 191, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b00100000; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10001101; c = 8'b10100001; // Expected: {'sum': 123, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10001101; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b00010001; c = 8'b00001101; // Expected: {'sum': 136, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b00010001; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01000010; c = 8'b00110011; // Expected: {'sum': 201, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01000010; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b11101110; c = 8'b11011000; // Expected: {'sum': 125, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b11101110; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11000100; c = 8'b10010000; // Expected: {'sum': 54, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11000100; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111001; b = 8'b11000011; c = 8'b10000110; // Expected: {'sum': 188, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111001; b = 8'b11000011; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b11010100; c = 8'b11100100; // Expected: {'sum': 81, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b11010100; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110100; c = 8'b01000000; // Expected: {'sum': 86, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110100; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11011101; c = 8'b11100100; // Expected: {'sum': 171, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11011101; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b10111001; c = 8'b01111000; // Expected: {'sum': 120, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b10111001; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10000111; c = 8'b11011001; // Expected: {'sum': 162, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10000111; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01001100; c = 8'b01101100; // Expected: {'sum': 106, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01001100; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 106, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10101001; c = 8'b00011111; // Expected: {'sum': 225, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10101001; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b00001000; c = 8'b01010000; // Expected: {'sum': 140, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b00001000; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11101101; c = 8'b10001100; // Expected: {'sum': 255, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11101101; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100001; b = 8'b00010111; c = 8'b01111111; // Expected: {'sum': 9, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100001; b = 8'b00010111; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b01100101; c = 8'b11110110; // Expected: {'sum': 203, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b01100101; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01001101; c = 8'b01101010; // Expected: {'sum': 48, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01001101; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b00000101; c = 8'b11100111; // Expected: {'sum': 176, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b00000101; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01110110; c = 8'b01100000; // Expected: {'sum': 161, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01110110; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01011110; c = 8'b00100011; // Expected: {'sum': 168, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01011110; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00010001; c = 8'b11000101; // Expected: {'sum': 144, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00010001; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00111011; c = 8'b11100100; // Expected: {'sum': 109, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00111011; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10010011; c = 8'b10110011; // Expected: {'sum': 75, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10010011; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b01110000; c = 8'b10010101; // Expected: {'sum': 48, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b01110000; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01111100; c = 8'b10001100; // Expected: {'sum': 33, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01111100; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111101; b = 8'b00001011; c = 8'b10100011; // Expected: {'sum': 85, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111101; b = 8'b00001011; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 85, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11100000; c = 8'b10010001; // Expected: {'sum': 68, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11100000; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b10010000; c = 8'b11100110; // Expected: {'sum': 177, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b10010000; c = 8'b11100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b01011000; c = 8'b10000110; // Expected: {'sum': 128, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b01011000; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b00001000; c = 8'b01101001; // Expected: {'sum': 30, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b00001000; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01000011; c = 8'b01110001; // Expected: {'sum': 154, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01000011; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b10101111; c = 8'b00101101; // Expected: {'sum': 121, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b10101111; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110100; b = 8'b11000011; c = 8'b01100010; // Expected: {'sum': 213, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110100; b = 8'b11000011; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b00111101; c = 8'b11100011; // Expected: {'sum': 209, 'carry': 47}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b00111101; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10010100; c = 8'b01111101; // Expected: {'sum': 13, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10010100; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b00001011; c = 8'b11000101; // Expected: {'sum': 154, 'carry': 69}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b00001011; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 154, 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00001100; c = 8'b00101000; // Expected: {'sum': 146, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00001100; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101000; b = 8'b10001001; c = 8'b01001000; // Expected: {'sum': 233, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101000; b = 8'b10001001; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000001; b = 8'b01111000; c = 8'b10110110; // Expected: {'sum': 143, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000001; b = 8'b01111000; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10101011; c = 8'b11100011; // Expected: {'sum': 94, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10101011; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11011011; c = 8'b11111110; // Expected: {'sum': 109, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11011011; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b01101111; c = 8'b11110100; // Expected: {'sum': 183, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b01101111; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b11011001; c = 8'b00011011; // Expected: {'sum': 56, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b11011001; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00111100; c = 8'b10011111; // Expected: {'sum': 199, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00111100; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b10101110; c = 8'b10011011; // Expected: {'sum': 68, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b10101110; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10111010; c = 8'b00100001; // Expected: {'sum': 2, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10111010; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b01101010; c = 8'b01010001; // Expected: {'sum': 74, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b01101010; c = 8'b01010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b10010111; c = 8'b01110000; // Expected: {'sum': 49, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b10010111; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b01000110; c = 8'b10110000; // Expected: {'sum': 51, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b01000110; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00001100; c = 8'b11100100; // Expected: {'sum': 81, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00001100; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11100111; c = 8'b10101100; // Expected: {'sum': 250, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11100111; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00100111; c = 8'b01001010; // Expected: {'sum': 65, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00100111; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00010010; c = 8'b01010101; // Expected: {'sum': 182, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00010010; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b00110000; c = 8'b00100100; // Expected: {'sum': 11, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b00110000; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2663,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11011110; c = 8'b00100101; // Expected: {'sum': 108, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11011110; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2664,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11101111; c = 8'b01111010; // Expected: {'sum': 129, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11101111; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2665,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01100111; c = 8'b00001001; // Expected: {'sum': 197, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01100111; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2666,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10010000; c = 8'b00001000; // Expected: {'sum': 112, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10010000; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2667,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b00001100; c = 8'b01010000; // Expected: {'sum': 80, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b00001100; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2668,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10001110; c = 8'b00001010; // Expected: {'sum': 0, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10001110; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2669,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00010011; c = 8'b01111001; // Expected: {'sum': 148, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00010011; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2670,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b00001000; c = 8'b11101101; // Expected: {'sum': 104, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b00001000; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2671,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b11110111; c = 8'b01011100; // Expected: {'sum': 59, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b11110111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2672,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11001001; c = 8'b00101110; // Expected: {'sum': 237, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11001001; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2673,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01110111; c = 8'b11111001; // Expected: {'sum': 71, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01110111; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2674,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b00010010; c = 8'b11011001; // Expected: {'sum': 190, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b00010010; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2675,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 190, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10010101; c = 8'b01010111; // Expected: {'sum': 148, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10010101; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2676,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10100010; c = 8'b11000010; // Expected: {'sum': 164, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10100010; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2677,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00001000; c = 8'b10000100; // Expected: {'sum': 62, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00001000; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2678,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01001110; c = 8'b01100101; // Expected: {'sum': 36, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01001110; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2679,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10110101; c = 8'b10111010; // Expected: {'sum': 201, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10110101; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2680,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11111001; c = 8'b10010001; // Expected: {'sum': 31, 'carry': 241}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11111001; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2681,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10011110; c = 8'b00100101; // Expected: {'sum': 8, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10011110; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2682,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10000110; c = 8'b10101111; // Expected: {'sum': 51, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10000110; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2683,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b11101111; c = 8'b00011101; // Expected: {'sum': 125, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b11101111; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2684,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b00010000; c = 8'b11100101; // Expected: {'sum': 228, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b00010000; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2685,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b10001100; c = 8'b00111100; // Expected: {'sum': 1, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b10001100; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2686,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b01010001; c = 8'b10010010; // Expected: {'sum': 54, 'carry': 209}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b01010001; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2687,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10100100; c = 8'b10010111; // Expected: {'sum': 86, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10100100; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2688,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00000101; c = 8'b00101101; // Expected: {'sum': 186, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00000101; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2689,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10111000; c = 8'b01000110; // Expected: {'sum': 239, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10111000; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2690,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11010011; c = 8'b11010110; // Expected: {'sum': 152, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11010011; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2691,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b01100011; c = 8'b11001100; // Expected: {'sum': 21, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b01100011; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2692,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100111; b = 8'b11010000; c = 8'b10111001; // Expected: {'sum': 78, 'carry': 177}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100111; b = 8'b11010000; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2693,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b00101001; c = 8'b00011011; // Expected: {'sum': 5, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b00101001; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2694,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b10000001; c = 8'b11101101; // Expected: {'sum': 18, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b10000001; c = 8'b11101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2695,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b00111110; c = 8'b10110100; // Expected: {'sum': 126, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b00111110; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2696,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b11011001; c = 8'b01101111; // Expected: {'sum': 6, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b11011001; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2697,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b11010000; c = 8'b10000101; // Expected: {'sum': 160, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b11010000; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2698,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10001101; c = 8'b01001101; // Expected: {'sum': 18, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10001101; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2699,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b10110100; c = 8'b00101000; // Expected: {'sum': 148, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b10110100; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2700,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b00110001; c = 8'b10101011; // Expected: {'sum': 197, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b00110001; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2701,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11111101; c = 8'b00110001; // Expected: {'sum': 216, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11111101; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2702,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11001011; c = 8'b01110010; // Expected: {'sum': 126, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11001011; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2703,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00110010; c = 8'b10010101; // Expected: {'sum': 26, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00110010; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2704,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b01100010; c = 8'b00001001; // Expected: {'sum': 197, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b01100010; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2705,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00101011; c = 8'b00011011; // Expected: {'sum': 28, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00101011; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2706,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b00011000; c = 8'b01111110; // Expected: {'sum': 32, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b00011000; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2707,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b01110111; c = 8'b10101101; // Expected: {'sum': 184, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b01110111; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2708,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b00100000; c = 8'b00011110; // Expected: {'sum': 36, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b00100000; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2709,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b10101110; c = 8'b11100001; // Expected: {'sum': 251, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b10101110; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2710,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b00101100; c = 8'b11100001; // Expected: {'sum': 240, 'carry': 45}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b00101100; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2711,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b01100010; c = 8'b10100001; // Expected: {'sum': 105, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b01100010; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2712,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b01100100; c = 8'b10111010; // Expected: {'sum': 36, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b01100100; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2713,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b10110010; c = 8'b11111001; // Expected: {'sum': 171, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b10110010; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2714,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11000111; c = 8'b01010011; // Expected: {'sum': 121, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11000111; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2715,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00001001; c = 8'b11100010; // Expected: {'sum': 202, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00001001; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2716,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11001000; c = 8'b10101110; // Expected: {'sum': 55, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11001000; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2717,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b10101110; c = 8'b10011000; // Expected: {'sum': 43, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b10101110; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2718,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01000010; c = 8'b01000111; // Expected: {'sum': 199, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01000010; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2719,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10111010; c = 8'b01010100; // Expected: {'sum': 176, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10111010; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2720,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00011110; c = 8'b01011010; // Expected: {'sum': 18, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00011110; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2721,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b00010101; c = 8'b11010001; // Expected: {'sum': 74, 'carry': 149}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b00010101; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2722,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10111000; c = 8'b01100111; // Expected: {'sum': 130, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10111000; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2723,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10100010; c = 8'b10100011; // Expected: {'sum': 47, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10100010; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2724,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b10010011; c = 8'b00100010; // Expected: {'sum': 233, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b10010011; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2725,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10111011; c = 8'b10000011; // Expected: {'sum': 22, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10111011; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2726,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 22, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11011001; c = 8'b10001100; // Expected: {'sum': 184, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11011001; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2727,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b01110010; c = 8'b01100111; // Expected: {'sum': 80, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b01110010; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2728,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 80, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01010111; c = 8'b10101010; // Expected: {'sum': 55, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01010111; c = 8'b10101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2729,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b01001111; c = 8'b11010001; // Expected: {'sum': 149, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b01001111; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2730,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10111010; c = 8'b01101011; // Expected: {'sum': 141, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10111010; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2731,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b10010011; c = 8'b00101001; // Expected: {'sum': 7, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b10010011; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2732,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b11000001; c = 8'b01011101; // Expected: {'sum': 90, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b11000001; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2733,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10111000; c = 8'b11100111; // Expected: {'sum': 217, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10111000; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2734,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10010110; c = 8'b00010001; // Expected: {'sum': 9, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10010110; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2735,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b10011000; c = 8'b01011111; // Expected: {'sum': 235, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b10011000; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2736,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b10011001; c = 8'b01111010; // Expected: {'sum': 116, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b10011001; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2737,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b11111010; c = 8'b00001011; // Expected: {'sum': 151, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b11111010; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2738,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10001101; c = 8'b11010000; // Expected: {'sum': 26, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10001101; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2739,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b01101000; c = 8'b11011111; // Expected: {'sum': 161, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b01101000; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2740,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10110100; c = 8'b00001101; // Expected: {'sum': 52, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10110100; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2741,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10011001; c = 8'b10001010; // Expected: {'sum': 54, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10011001; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2742,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001111; b = 8'b01101000; c = 8'b11001000; // Expected: {'sum': 111, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001111; b = 8'b01101000; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2743,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b11010111; c = 8'b00101100; // Expected: {'sum': 23, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b11010111; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2744,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10011010; c = 8'b01011110; // Expected: {'sum': 243, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10011010; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2745,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11100111; c = 8'b00000100; // Expected: {'sum': 95, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11100111; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2746,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b10011010; c = 8'b01101100; // Expected: {'sum': 91, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b10011010; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2747,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10111000; c = 8'b01101010; // Expected: {'sum': 58, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10111000; c = 8'b01101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2748,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00100101; c = 8'b11000100; // Expected: {'sum': 74, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00100101; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2749,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b10001111; c = 8'b01010101; // Expected: {'sum': 145, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b10001111; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2750,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11100010; c = 8'b11011010; // Expected: {'sum': 102, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11100010; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2751,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01101000; c = 8'b01101001; // Expected: {'sum': 75, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01101000; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2752,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01011001; c = 8'b11011101; // Expected: {'sum': 209, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01011001; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2753,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b00101010; c = 8'b10101001; // Expected: {'sum': 100, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b00101010; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2754,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b11101011; c = 8'b00111100; // Expected: {'sum': 40, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b11101011; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2755,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b01001010; c = 8'b11111111; // Expected: {'sum': 88, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b01001010; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2756,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00010001; c = 8'b11001011; // Expected: {'sum': 249, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00010001; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2757,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b00111101; c = 8'b10011101; // Expected: {'sum': 12, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b00111101; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2758,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00010011; c = 8'b10001111; // Expected: {'sum': 143, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00010011; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2759,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b01001011; c = 8'b00100010; // Expected: {'sum': 173, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b01001011; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2760,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01110000; c = 8'b01000110; // Expected: {'sum': 105, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01110000; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2761,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10111010; c = 8'b10010011; // Expected: {'sum': 58, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10111010; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2762,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01110000; c = 8'b11010011; // Expected: {'sum': 92, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01110000; c = 8'b11010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2763,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00011111; c = 8'b11100111; // Expected: {'sum': 69, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00011111; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2764,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00011110; c = 8'b01001011; // Expected: {'sum': 143, 'carry': 90}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00011110; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2765,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b01000010; c = 8'b11101110; // Expected: {'sum': 83, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b01000010; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2766,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01011100; c = 8'b00111010; // Expected: {'sum': 123, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01011100; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2767,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10110000; c = 8'b01011000; // Expected: {'sum': 228, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10110000; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2768,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b11001011; c = 8'b01001001; // Expected: {'sum': 185, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b11001011; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2769,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b01111000; c = 8'b00011010; // Expected: {'sum': 8, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b01111000; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2770,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b11110110; c = 8'b10011110; // Expected: {'sum': 205, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b11110110; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2771,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10001100; c = 8'b10010111; // Expected: {'sum': 211, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10001100; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2772,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10011011; c = 8'b00001000; // Expected: {'sum': 227, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10011011; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2773,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b01001111; c = 8'b10011011; // Expected: {'sum': 68, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b01001111; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2774,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b11010001; c = 8'b11011110; // Expected: {'sum': 185, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b11010001; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2775,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b10111100; c = 8'b11000100; // Expected: {'sum': 103, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b10111100; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2776,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11110111; c = 8'b10111001; // Expected: {'sum': 60, 'carry': 243}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11110111; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2777,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11000111; c = 8'b01100010; // Expected: {'sum': 128, 'carry': 103}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11000111; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2778,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100010; b = 8'b11111011; c = 8'b10000011; // Expected: {'sum': 90, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100010; b = 8'b11111011; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2779,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b00101100; c = 8'b01111110; // Expected: {'sum': 120, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b00101100; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2780,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b00011010; c = 8'b10000111; // Expected: {'sum': 48, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b00011010; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2781,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b11110110; c = 8'b11110110; // Expected: {'sum': 130, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b11110110; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2782,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11000010; c = 8'b01111101; // Expected: {'sum': 137, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11000010; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2783,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10001010; c = 8'b00100101; // Expected: {'sum': 94, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10001010; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2784,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b01110110; c = 8'b11100010; // Expected: {'sum': 221, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b01110110; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2785,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b11100110; c = 8'b10000100; // Expected: {'sum': 193, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b11100110; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2786,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011010; b = 8'b00001101; c = 8'b00010100; // Expected: {'sum': 195, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011010; b = 8'b00001101; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2787,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00110111; c = 8'b01110000; // Expected: {'sum': 107, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00110111; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2788,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b11000010; c = 8'b11001010; // Expected: {'sum': 9, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b11000010; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2789,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00011111; c = 8'b01010110; // Expected: {'sum': 215, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00011111; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2790,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10011101; c = 8'b00100110; // Expected: {'sum': 20, 'carry': 175}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10011101; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2791,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10111110; c = 8'b00101110; // Expected: {'sum': 66, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10111110; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2792,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b11111010; c = 8'b01101110; // Expected: {'sum': 170, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b11111010; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2793,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01110001; c = 8'b10001110; // Expected: {'sum': 4, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01110001; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2794,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11010111; c = 8'b10100010; // Expected: {'sum': 226, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11010111; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2795,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11100011; c = 8'b00101011; // Expected: {'sum': 41, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11100011; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2796,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b10111001; c = 8'b00110000; // Expected: {'sum': 136, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b10111001; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2797,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10100001; c = 8'b01100011; // Expected: {'sum': 89, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10100001; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2798,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b01111010; c = 8'b11110111; // Expected: {'sum': 34, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b01111010; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2799,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b10010011; c = 8'b01010011; // Expected: {'sum': 128, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b10010011; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2800,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b00101100; c = 8'b00001001; // Expected: {'sum': 213, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b00101100; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2801,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b01011110; c = 8'b10011010; // Expected: {'sum': 56, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b01011110; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2802,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b01111010; c = 8'b00000110; // Expected: {'sum': 238, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b01111010; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2803,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b11100111; c = 8'b00110001; // Expected: {'sum': 82, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b11100111; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2804,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b01011000; c = 8'b11011010; // Expected: {'sum': 93, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b01011000; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2805,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b00101010; c = 8'b01001000; // Expected: {'sum': 147, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b00101010; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2806,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b11101011; c = 8'b10101001; // Expected: {'sum': 220, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b11101011; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2807,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b00111011; c = 8'b11001011; // Expected: {'sum': 218, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b00111011; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2808,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00001011; c = 8'b11000000; // Expected: {'sum': 73, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00001011; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2809,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01001110; c = 8'b11001011; // Expected: {'sum': 58, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01001110; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2810,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10010100; c = 8'b00110110; // Expected: {'sum': 4, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10010100; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2811,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b11001101; c = 8'b11010101; // Expected: {'sum': 66, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b11001101; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2812,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b11011010; c = 8'b01100010; // Expected: {'sum': 42, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b11011010; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2813,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b11010101; c = 8'b00010010; // Expected: {'sum': 250, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b11010101; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2814,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010001; b = 8'b01100101; c = 8'b01101110; // Expected: {'sum': 218, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010001; b = 8'b01100101; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2815,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b00010000; c = 8'b10111100; // Expected: {'sum': 234, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b00010000; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2816,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010000; b = 8'b10110110; c = 8'b00000100; // Expected: {'sum': 34, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010000; b = 8'b10110110; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2817,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10011111; c = 8'b01101011; // Expected: {'sum': 226, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10011111; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2818,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10111111; c = 8'b00111010; // Expected: {'sum': 29, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10111111; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2819,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b11111101; c = 8'b10111110; // Expected: {'sum': 196, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b11111101; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2820,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11111001; c = 8'b11010101; // Expected: {'sum': 187, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11111001; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2821,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10101111; c = 8'b11111110; // Expected: {'sum': 230, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10101111; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2822,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10000010; c = 8'b00000101; // Expected: {'sum': 68, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10000010; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2823,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b01010001; c = 8'b11001011; // Expected: {'sum': 26, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b01010001; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2824,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b01001101; c = 8'b11001110; // Expected: {'sum': 13, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b01001101; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2825,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11101001; c = 8'b00000100; // Expected: {'sum': 9, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11101001; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2826,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100111; b = 8'b11011111; c = 8'b00110000; // Expected: {'sum': 72, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100111; b = 8'b11011111; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2827,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b11000110; c = 8'b11001011; // Expected: {'sum': 55, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b11000110; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2828,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b11001000; c = 8'b00001001; // Expected: {'sum': 136, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b11001000; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2829,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000101; b = 8'b00011110; c = 8'b00101011; // Expected: {'sum': 48, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000101; b = 8'b00011110; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2830,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b00001010; c = 8'b11111001; // Expected: {'sum': 214, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b00001010; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2831,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b00111011; c = 8'b11000111; // Expected: {'sum': 68, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b00111011; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2832,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10011111; c = 8'b11101011; // Expected: {'sum': 224, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10011111; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2833,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10011110; c = 8'b11001110; // Expected: {'sum': 227, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10011110; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2834,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b11000111; c = 8'b00100000; // Expected: {'sum': 91, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b11000111; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2835,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b11101010; c = 8'b10011011; // Expected: {'sum': 87, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b11101010; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2836,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01001011; c = 8'b00010100; // Expected: {'sum': 39, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01001011; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2837,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10110000; c = 8'b10010000; // Expected: {'sum': 245, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10110000; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2838,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b01010110; c = 8'b10101001; // Expected: {'sum': 223, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b01010110; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2839,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b01110100; c = 8'b00011011; // Expected: {'sum': 206, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b01110100; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2840,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01010101; c = 8'b11001110; // Expected: {'sum': 145, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01010101; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2841,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b11011010; c = 8'b10010111; // Expected: {'sum': 99, 'carry': 158}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b11011010; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2842,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10101000; c = 8'b11001011; // Expected: {'sum': 50, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10101000; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2843,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11100110; c = 8'b01010011; // Expected: {'sum': 36, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11100110; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2844,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11010110; c = 8'b10111101; // Expected: {'sum': 139, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11010110; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2845,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b01000000; c = 8'b00100000; // Expected: {'sum': 57, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b01000000; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2846,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b00100111; c = 8'b10010101; // Expected: {'sum': 122, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b00100111; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2847,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11010000; c = 8'b00010101; // Expected: {'sum': 223, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11010000; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2848,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b10010011; c = 8'b00101100; // Expected: {'sum': 128, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b10010011; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2849,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b11101001; c = 8'b10100011; // Expected: {'sum': 117, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b11101001; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2850,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 117, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b11110001; c = 8'b10001011; // Expected: {'sum': 212, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b11110001; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2851,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b11001011; c = 8'b00001100; // Expected: {'sum': 187, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b11001011; c = 8'b00001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2852,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b10011111; c = 8'b01111000; // Expected: {'sum': 212, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b10011111; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2853,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00000111; c = 8'b10000011; // Expected: {'sum': 26, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00000111; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2854,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b10001100; c = 8'b11010000; // Expected: {'sum': 158, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b10001100; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2855,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b10101110; c = 8'b01111100; // Expected: {'sum': 219, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b10101110; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2856,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b11000101; c = 8'b01011010; // Expected: {'sum': 104, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b11000101; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2857,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b01010000; c = 8'b10000111; // Expected: {'sum': 192, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b01010000; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2858,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b01111010; c = 8'b11001111; // Expected: {'sum': 14, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b01111010; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2859,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b10111101; c = 8'b01001111; // Expected: {'sum': 166, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b10111101; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2860,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00000100; c = 8'b11101011; // Expected: {'sum': 175, 'carry': 64}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00000100; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2861,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10011001; c = 8'b01111101; // Expected: {'sum': 217, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10011001; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2862,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b10111001; c = 8'b10011101; // Expected: {'sum': 81, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b10111001; c = 8'b10011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2863,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b00011010; c = 8'b10011011; // Expected: {'sum': 35, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b00011010; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2864,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011100; b = 8'b00001111; c = 8'b11000111; // Expected: {'sum': 212, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011100; b = 8'b00001111; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2865,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b00101111; c = 8'b11000011; // Expected: {'sum': 10, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b00101111; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2866,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b00110101; c = 8'b00101011; // Expected: {'sum': 61, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b00110101; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2867,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00011100; c = 8'b11011110; // Expected: {'sum': 98, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00011100; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2868,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b01111100; c = 8'b11011000; // Expected: {'sum': 130, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b01111100; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2869,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b01100011; c = 8'b00011001; // Expected: {'sum': 220, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b01100011; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2870,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b00000110; c = 8'b01010000; // Expected: {'sum': 43, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b00000110; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2871,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11100110; c = 8'b01111000; // Expected: {'sum': 162, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11100110; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2872,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01010011; c = 8'b00100100; // Expected: {'sum': 175, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01010011; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2873,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b01000101; c = 8'b10000010; // Expected: {'sum': 120, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b01000101; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2874,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01000010; c = 8'b00011100; // Expected: {'sum': 176, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01000010; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2875,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 176, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11110011; c = 8'b11100111; // Expected: {'sum': 29, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11110011; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2876,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b10110000; c = 8'b11101111; // Expected: {'sum': 228, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b10110000; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2877,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01011111; c = 8'b10101100; // Expected: {'sum': 174, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01011111; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2878,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00001001; c = 8'b10111100; // Expected: {'sum': 20, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00001001; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2879,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b11110000; c = 8'b00011101; // Expected: {'sum': 247, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b11110000; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2880,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b01011011; c = 8'b10000010; // Expected: {'sum': 226, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b01011011; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2881,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00110101; c = 8'b11100011; // Expected: {'sum': 214, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00110101; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2882,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b10010100; c = 8'b10000000; // Expected: {'sum': 75, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b10010100; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2883,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00101001; c = 8'b01111110; // Expected: {'sum': 20, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00101001; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2884,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b01110000; c = 8'b01000010; // Expected: {'sum': 172, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b01110000; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2885,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b11100100; c = 8'b01001100; // Expected: {'sum': 136, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b11100100; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2886,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10010011; c = 8'b00010110; // Expected: {'sum': 207, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10010011; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2887,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b00000010; c = 8'b10010000; // Expected: {'sum': 152, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b00000010; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2888,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10011111; c = 8'b10100101; // Expected: {'sum': 82, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10011111; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2889,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000011; b = 8'b11000101; c = 8'b01110010; // Expected: {'sum': 180, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000011; b = 8'b11000101; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2890,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b00101000; c = 8'b00101011; // Expected: {'sum': 47, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b00101000; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2891,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b01000100; c = 8'b11110101; // Expected: {'sum': 2, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b01000100; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2892,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11011101; c = 8'b00100101; // Expected: {'sum': 238, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11011101; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2893,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 238, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b00101000; c = 8'b01101111; // Expected: {'sum': 16, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b00101000; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2894,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01010100; c = 8'b11100011; // Expected: {'sum': 219, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01010100; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2895,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b11101110; c = 8'b00001011; // Expected: {'sum': 15, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b11101110; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2896,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b01111001; c = 8'b00001010; // Expected: {'sum': 40, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b01111001; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2897,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b00000100; c = 8'b01001100; // Expected: {'sum': 200, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b00000100; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2898,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00010010; c = 8'b00111011; // Expected: {'sum': 254, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00010010; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2899,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b10111111; c = 8'b10010100; // Expected: {'sum': 2, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b10111111; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2900,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b00111100; c = 8'b10000000; // Expected: {'sum': 180, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b00111100; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2901,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b10001101; c = 8'b00111101; // Expected: {'sum': 21, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b10001101; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2902,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b11011110; c = 8'b00101010; // Expected: {'sum': 157, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b11011110; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2903,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10000110; c = 8'b00011100; // Expected: {'sum': 87, 'carry': 140}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10000110; c = 8'b00011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2904,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 87, 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b01000110; c = 8'b01000001; // Expected: {'sum': 113, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b01000110; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2905,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b01100001; c = 8'b00011011; // Expected: {'sum': 125, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b01100001; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2906,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b10101111; c = 8'b01000111; // Expected: {'sum': 112, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b10101111; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2907,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b01011100; c = 8'b01000011; // Expected: {'sum': 217, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b01011100; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2908,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b11100100; c = 8'b00111100; // Expected: {'sum': 60, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b11100100; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2909,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b11100101; c = 8'b00111111; // Expected: {'sum': 216, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b11100101; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2910,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10100100; c = 8'b00001101; // Expected: {'sum': 236, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10100100; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2911,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b11011111; c = 8'b00110001; // Expected: {'sum': 187, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b11011111; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2912,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b10100101; c = 8'b00010101; // Expected: {'sum': 50, 'carry': 133}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b10100101; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2913,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b01000111; c = 8'b11010000; // Expected: {'sum': 81, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b01000111; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2914,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 81, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11010110; c = 8'b00000111; // Expected: {'sum': 101, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11010110; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2915,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b00010110; c = 8'b11101000; // Expected: {'sum': 104, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b00010110; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2916,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00110000; c = 8'b01011001; // Expected: {'sum': 183, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00110000; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2917,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b11011111; c = 8'b01101011; // Expected: {'sum': 157, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b11011111; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2918,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b00010110; c = 8'b00100101; // Expected: {'sum': 118, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b00010110; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2919,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01000011; c = 8'b01011100; // Expected: {'sum': 140, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01000011; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2920,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00111001; c = 8'b01111011; // Expected: {'sum': 241, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00111001; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2921,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110001; b = 8'b00111011; c = 8'b01010100; // Expected: {'sum': 94, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110001; b = 8'b00111011; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2922,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b01000110; c = 8'b10001101; // Expected: {'sum': 251, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b01000110; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2923,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11110010; c = 8'b11001100; // Expected: {'sum': 175, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11110010; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2924,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b11010010; c = 8'b00011000; // Expected: {'sum': 218, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b11010010; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2925,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11111101; c = 8'b01100011; // Expected: {'sum': 58, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11111101; c = 8'b01100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2926,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b10111100; c = 8'b00110010; // Expected: {'sum': 245, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b10111100; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2927,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b10110111; c = 8'b10111000; // Expected: {'sum': 50, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b10110111; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2928,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b11010001; c = 8'b10000110; // Expected: {'sum': 215, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b11010001; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2929,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b01010111; c = 8'b00010110; // Expected: {'sum': 170, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b01010111; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2930,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b11110010; c = 8'b10110100; // Expected: {'sum': 135, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b11110010; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2931,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b01010110; c = 8'b01100110; // Expected: {'sum': 227, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b01010110; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2932,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b10010100; c = 8'b01001110; // Expected: {'sum': 157, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b10010100; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2933,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10111000; c = 8'b11011010; // Expected: {'sum': 218, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10111000; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2934,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b00001101; c = 8'b10100101; // Expected: {'sum': 102, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b00001101; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2935,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 102, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10111101; c = 8'b00010100; // Expected: {'sum': 15, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10111101; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2936,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b00000111; c = 8'b01110101; // Expected: {'sum': 1, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b00000111; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2937,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11101011; c = 8'b01000110; // Expected: {'sum': 53, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11101011; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2938,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00101001; c = 8'b01101001; // Expected: {'sum': 57, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00101001; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2939,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10111110; c = 8'b10101111; // Expected: {'sum': 206, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10111110; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2940,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10100000; c = 8'b01110000; // Expected: {'sum': 198, 'carry': 48}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10100000; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2941,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10011111; c = 8'b10100100; // Expected: {'sum': 35, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10011111; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2942,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01100101; c = 8'b10100001; // Expected: {'sum': 120, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01100101; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2943,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b10011101; c = 8'b10010011; // Expected: {'sum': 112, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b10011101; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2944,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00000010; c = 8'b01101000; // Expected: {'sum': 14, 'carry': 96}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00000010; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2945,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10111110; c = 8'b00110000; // Expected: {'sum': 137, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10111110; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2946,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010011; b = 8'b01110010; c = 8'b00111111; // Expected: {'sum': 30, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010011; b = 8'b01110010; c = 8'b00111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2947,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b01111111; c = 8'b11100000; // Expected: {'sum': 179, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b01111111; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2948,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01010010; c = 8'b00101011; // Expected: {'sum': 121, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01010010; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2949,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b01011100; c = 8'b00011101; // Expected: {'sum': 214, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b01011100; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2950,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00001010; c = 8'b01010100; // Expected: {'sum': 29, 'carry': 66}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00001010; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2951,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10000011; c = 8'b10100111; // Expected: {'sum': 65, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10000011; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2952,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10100111; c = 8'b11010101; // Expected: {'sum': 64, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10100111; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2953,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01011101; c = 8'b00111001; // Expected: {'sum': 107, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01011101; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2954,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 107, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b00011000; c = 8'b11100011; // Expected: {'sum': 163, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b00011000; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2955,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111010; b = 8'b00110100; c = 8'b01001110; // Expected: {'sum': 0, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111010; b = 8'b00110100; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2956,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01100111; c = 8'b00110001; // Expected: {'sum': 179, 'carry': 101}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01100111; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2957,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b01101110; c = 8'b11110010; // Expected: {'sum': 168, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b01101110; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2958,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11101000; c = 8'b01010000; // Expected: {'sum': 41, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11101000; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2959,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b10000100; c = 8'b00000011; // Expected: {'sum': 178, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b10000100; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2960,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b11101111; c = 8'b00101010; // Expected: {'sum': 71, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b11101111; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2961,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00000001; c = 8'b00101000; // Expected: {'sum': 116, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00000001; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2962,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11101001; c = 8'b01010100; // Expected: {'sum': 98, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11101001; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2963,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b10101110; c = 8'b01101000; // Expected: {'sum': 91, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b10101110; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2964,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 91, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b01010010; c = 8'b10100101; // Expected: {'sum': 251, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b01010010; c = 8'b10100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2965,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01100111; c = 8'b10101011; // Expected: {'sum': 71, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01100111; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2966,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000010; b = 8'b00010101; c = 8'b10101000; // Expected: {'sum': 63, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000010; b = 8'b00010101; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2967,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b00010101; c = 8'b00011101; // Expected: {'sum': 208, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b00010101; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2968,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00011110; c = 8'b11011110; // Expected: {'sum': 30, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00011110; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2969,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10100101; c = 8'b01111100; // Expected: {'sum': 29, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10100101; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2970,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b11111101; c = 8'b10100001; // Expected: {'sum': 248, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b11111101; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2971,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11111111; c = 8'b01101001; // Expected: {'sum': 68, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11111111; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2972,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b11001011; c = 8'b00100001; // Expected: {'sum': 221, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b11001011; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2973,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b11111010; c = 8'b11001100; // Expected: {'sum': 199, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b11111010; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2974,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b10110011; c = 8'b00000110; // Expected: {'sum': 94, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b10110011; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2975,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b11101011; c = 8'b00110100; // Expected: {'sum': 216, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b11101011; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2976,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b11110001; c = 8'b00111000; // Expected: {'sum': 151, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b11110001; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2977,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00011100; c = 8'b11110010; // Expected: {'sum': 92, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00011100; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2978,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b00010101; c = 8'b01001001; // Expected: {'sum': 143, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b00010101; c = 8'b01001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2979,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00110001; c = 8'b10111001; // Expected: {'sum': 119, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00110001; c = 8'b10111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2980,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01100110; c = 8'b10000111; // Expected: {'sum': 171, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01100110; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2981,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b10011100; c = 8'b00100110; // Expected: {'sum': 95, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b10011100; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2982,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b11111100; c = 8'b11000111; // Expected: {'sum': 46, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b11111100; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2983,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b01011111; c = 8'b00110110; // Expected: {'sum': 125, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b01011111; c = 8'b00110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2984,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11101001; c = 8'b00011110; // Expected: {'sum': 130, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11101001; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2985,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01100001; c = 8'b11000011; // Expected: {'sum': 62, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01100001; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2986,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11100111; c = 8'b10101011; // Expected: {'sum': 139, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11100111; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2987,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b00100000; c = 8'b10101111; // Expected: {'sum': 182, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b00100000; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2988,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001110; b = 8'b00111010; c = 8'b10101011; // Expected: {'sum': 223, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001110; b = 8'b00111010; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2989,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b01011001; c = 8'b11111000; // Expected: {'sum': 147, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b01011001; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2990,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b01010100; c = 8'b10110110; // Expected: {'sum': 103, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b01010100; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2991,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10001010; c = 8'b11010100; // Expected: {'sum': 92, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10001010; c = 8'b11010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2992,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b11001011; c = 8'b00111110; // Expected: {'sum': 230, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b11001011; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2993,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00100011; c = 8'b11000111; // Expected: {'sum': 98, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00100011; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2994,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b00101000; c = 8'b00101111; // Expected: {'sum': 196, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b00101000; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2995,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11001111; c = 8'b01111111; // Expected: {'sum': 149, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11001111; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2996,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10000100; c = 8'b10101110; // Expected: {'sum': 124, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10000100; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2997,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 124, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01011001; c = 8'b11011011; // Expected: {'sum': 90, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01011001; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2998,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010010; b = 8'b10010100; c = 8'b11100000; // Expected: {'sum': 38, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010010; b = 8'b10010100; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2999,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b00001100; c = 8'b00101101; // Expected: {'sum': 47, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b00001100; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3000,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b01100010; c = 8'b00100000; // Expected: {'sum': 222, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b01100010; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3001,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b10001011; c = 8'b10101000; // Expected: {'sum': 146, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b10001011; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3002,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b01001011; c = 8'b00101100; // Expected: {'sum': 40, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b01001011; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3003,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b00001100; c = 8'b00110100; // Expected: {'sum': 179, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b00001100; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3004,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00010100; c = 8'b00110100; // Expected: {'sum': 222, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00010100; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3005,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b11100101; c = 8'b10101000; // Expected: {'sum': 193, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b11100101; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3006,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10011010; c = 8'b01001011; // Expected: {'sum': 29, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10011010; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3007,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b11001000; c = 8'b01101100; // Expected: {'sum': 213, 'carry': 104}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b11001000; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3008,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11000100; c = 8'b11010010; // Expected: {'sum': 51, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11000100; c = 8'b11010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3009,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b00000011; c = 8'b11101100; // Expected: {'sum': 82, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b00000011; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3010,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b11010101; c = 8'b01100001; // Expected: {'sum': 254, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b11010101; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3011,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b10010111; c = 8'b11001000; // Expected: {'sum': 58, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b10010111; c = 8'b11001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3012,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b01111110; c = 8'b01110110; // Expected: {'sum': 125, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b01111110; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3013,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01111101; c = 8'b00000110; // Expected: {'sum': 46, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01111101; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3014,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b10011001; c = 8'b10101111; // Expected: {'sum': 92, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b10011001; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3015,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b00000111; c = 8'b01111001; // Expected: {'sum': 21, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b00000111; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3016,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b01100101; c = 8'b10000110; // Expected: {'sum': 172, 'carry': 71}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b01100101; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3017,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11010110; c = 8'b01111110; // Expected: {'sum': 255, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11010110; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3018,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b01101100; c = 8'b00011101; // Expected: {'sum': 13, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b01101100; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3019,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b11011000; c = 8'b00010111; // Expected: {'sum': 188, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b11011000; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3020,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b11001011; c = 8'b11110110; // Expected: {'sum': 67, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b11001011; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3021,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b10001010; c = 8'b00110111; // Expected: {'sum': 49, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b10001010; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3022,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b10000001; c = 8'b00000110; // Expected: {'sum': 164, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b10000001; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3023,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00011011; c = 8'b11011001; // Expected: {'sum': 23, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00011011; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3024,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b10011000; c = 8'b10011111; // Expected: {'sum': 67, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b10011000; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3025,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b01001000; c = 8'b00111011; // Expected: {'sum': 160, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b01001000; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3026,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11100100; c = 8'b11000011; // Expected: {'sum': 245, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11100100; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3027,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b11111000; c = 8'b01001010; // Expected: {'sum': 110, 'carry': 216}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b11111000; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3028,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11111100; c = 8'b11001001; // Expected: {'sum': 100, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11111100; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3029,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10000011; c = 8'b10000111; // Expected: {'sum': 65, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10000011; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3030,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b10100011; c = 8'b10000010; // Expected: {'sum': 63, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b10100011; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3031,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01011001; c = 8'b00001010; // Expected: {'sum': 148, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01011001; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3032,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11000000; c = 8'b11100100; // Expected: {'sum': 228, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11000000; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3033,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b01001110; c = 8'b11110010; // Expected: {'sum': 8, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b01001110; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3034,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10010111; c = 8'b00100011; // Expected: {'sum': 31, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10010111; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3035,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b10000101; c = 8'b00001011; // Expected: {'sum': 31, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b10000101; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3036,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10101111; c = 8'b00010000; // Expected: {'sum': 119, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10101111; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3037,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b10110111; c = 8'b11110111; // Expected: {'sum': 23, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b10110111; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3038,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b01101011; c = 8'b11001001; // Expected: {'sum': 14, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b01101011; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3039,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b11100111; c = 8'b01001000; // Expected: {'sum': 120, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b11100111; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3040,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b10010000; c = 8'b00011000; // Expected: {'sum': 76, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b10010000; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3041,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10111001; c = 8'b10111000; // Expected: {'sum': 3, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10111001; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3042,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b10000111; c = 8'b10000011; // Expected: {'sum': 224, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b10000111; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3043,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b00000100; c = 8'b00100110; // Expected: {'sum': 185, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b00000100; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3044,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b10111110; c = 8'b00011101; // Expected: {'sum': 243, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b10111110; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3045,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b11100001; c = 8'b10001110; // Expected: {'sum': 104, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b11100001; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3046,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b10101010; c = 8'b01000001; // Expected: {'sum': 128, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b10101010; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3047,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11100001; c = 8'b10111111; // Expected: {'sum': 86, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11100001; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3048,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b01110111; c = 8'b01010110; // Expected: {'sum': 232, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b01110111; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3049,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b11000011; c = 8'b01100101; // Expected: {'sum': 75, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b11000011; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3050,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11111100; c = 8'b11100100; // Expected: {'sum': 169, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11111100; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3051,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b01100100; c = 8'b00100011; // Expected: {'sum': 254, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b01100100; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3052,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b00000100; c = 8'b00000111; // Expected: {'sum': 153, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b00000100; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3053,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b00100000; c = 8'b01001010; // Expected: {'sum': 233, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b00100000; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3054,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01011100; c = 8'b00001010; // Expected: {'sum': 41, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01011100; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3055,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b01011100; c = 8'b10001010; // Expected: {'sum': 1, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b01011100; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3056,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10111010; c = 8'b01101101; // Expected: {'sum': 196, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10111010; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3057,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00100100; c = 8'b01001101; // Expected: {'sum': 38, 'carry': 77}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00100100; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3058,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b00111101; c = 8'b11101011; // Expected: {'sum': 195, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b00111101; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3059,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 195, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b10010011; c = 8'b10010110; // Expected: {'sum': 210, 'carry': 151}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b10010011; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3060,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11110001; c = 8'b10100111; // Expected: {'sum': 43, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11110001; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3061,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 43, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b11001111; c = 8'b01011100; // Expected: {'sum': 148, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b11001111; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3062,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00110011; c = 8'b10000111; // Expected: {'sum': 153, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00110011; c = 8'b10000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3063,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10110111; c = 8'b00001000; // Expected: {'sum': 225, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10110111; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3064,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11010100; c = 8'b00101001; // Expected: {'sum': 209, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11010100; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3065,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b10001001; c = 8'b10110110; // Expected: {'sum': 88, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b10001001; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3066,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 88, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11011000; c = 8'b11010001; // Expected: {'sum': 48, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11011000; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3067,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b00001100; c = 8'b01011111; // Expected: {'sum': 203, 'carry': 28}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b00001100; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3068,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b01110001; c = 8'b11011100; // Expected: {'sum': 148, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b01110001; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3069,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b11000010; c = 8'b10010010; // Expected: {'sum': 112, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b11000010; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3070,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b10010111; c = 8'b11100111; // Expected: {'sum': 126, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b10010111; c = 8'b11100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3071,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b11100101; c = 8'b10101001; // Expected: {'sum': 241, 'carry': 173}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b11100101; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3072,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001011; b = 8'b01100111; c = 8'b00110111; // Expected: {'sum': 219, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001011; b = 8'b01100111; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3073,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01001010; c = 8'b00111110; // Expected: {'sum': 149, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01001010; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3074,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011001; b = 8'b10111011; c = 8'b11001111; // Expected: {'sum': 173, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011001; b = 8'b10111011; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3075,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000011; b = 8'b01001110; c = 8'b01011101; // Expected: {'sum': 144, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000011; b = 8'b01001110; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3076,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 144, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b10101000; c = 8'b10100011; // Expected: {'sum': 9, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b10101000; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3077,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101111; b = 8'b00000111; c = 8'b00011011; // Expected: {'sum': 51, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101111; b = 8'b00000111; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3078,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b11101100; c = 8'b00101010; // Expected: {'sum': 32, 'carry': 238}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b11101100; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3079,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 32, 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10010010; c = 8'b01101111; // Expected: {'sum': 232, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10010010; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3080,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01110001; c = 8'b00000001; // Expected: {'sum': 246, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01110001; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3081,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 246, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b10010100; c = 8'b01111011; // Expected: {'sum': 35, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b10010100; c = 8'b01111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3082,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10110000; c = 8'b11000010; // Expected: {'sum': 131, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10110000; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3083,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b11111111; c = 8'b00000100; // Expected: {'sum': 83, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b11111111; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3084,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b01011011; c = 8'b11000010; // Expected: {'sum': 126, 'carry': 195}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b01011011; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3085,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10000101; c = 8'b11101010; // Expected: {'sum': 104, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10000101; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3086,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10110111; c = 8'b00111010; // Expected: {'sum': 129, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10110111; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3087,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10110110; c = 8'b11100011; // Expected: {'sum': 162, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10110110; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3088,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b10011101; c = 8'b01001111; // Expected: {'sum': 229, 'carry': 31}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b10011101; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3089,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 229, 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b10001110; c = 8'b10000110; // Expected: {'sum': 224, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b10001110; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3090,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b11001010; c = 8'b00011111; // Expected: {'sum': 196, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b11001010; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3091,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001101; b = 8'b10100000; c = 8'b10101100; // Expected: {'sum': 193, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001101; b = 8'b10100000; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3092,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b01111010; c = 8'b00100001; // Expected: {'sum': 10, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b01111010; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3093,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b10100000; c = 8'b00010100; // Expected: {'sum': 159, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b10100000; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3094,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11010111; c = 8'b00111010; // Expected: {'sum': 180, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11010111; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3095,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10000011; c = 8'b00011011; // Expected: {'sum': 141, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10000011; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3096,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01011101; c = 8'b10111100; // Expected: {'sum': 104, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01011101; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3097,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 104, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b00111101; c = 8'b00010000; // Expected: {'sum': 253, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b00111101; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3098,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b10100111; c = 8'b01110010; // Expected: {'sum': 66, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b10100111; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3099,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10101111; c = 8'b00011001; // Expected: {'sum': 95, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10101111; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00100010; c = 8'b01111110; // Expected: {'sum': 239, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00100010; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10001010; c = 8'b00100000; // Expected: {'sum': 210, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10001010; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01100111; c = 8'b01010011; // Expected: {'sum': 159, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01100111; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b01011000; c = 8'b11101110; // Expected: {'sum': 78, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b01011000; c = 8'b11101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b11110111; c = 8'b00001110; // Expected: {'sum': 71, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b11110111; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b10110011; c = 8'b01000000; // Expected: {'sum': 232, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b10110011; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01001111; c = 8'b00100111; // Expected: {'sum': 7, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01001111; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11000010; c = 8'b10011100; // Expected: {'sum': 9, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11000010; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b00111100; c = 8'b10111101; // Expected: {'sum': 7, 'carry': 188}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b00111100; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b11110100; c = 8'b00100011; // Expected: {'sum': 8, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b11110100; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b00111000; c = 8'b11111001; // Expected: {'sum': 105, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b00111000; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b10001101; c = 8'b00010110; // Expected: {'sum': 114, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b10001101; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00010011; c = 8'b00010010; // Expected: {'sum': 179, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00010011; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b10010111; c = 8'b11111111; // Expected: {'sum': 208, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b10010111; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b11011000; c = 8'b00010001; // Expected: {'sum': 94, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b11011000; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b11011000; c = 8'b10010000; // Expected: {'sum': 120, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b11011000; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10100111; c = 8'b11001001; // Expected: {'sum': 159, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10100111; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10100001; c = 8'b00000001; // Expected: {'sum': 6, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10100001; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10100000; c = 8'b00000001; // Expected: {'sum': 185, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10100000; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11110000; c = 8'b11110000; // Expected: {'sum': 30, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11110000; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b11100101; c = 8'b11011001; // Expected: {'sum': 58, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b11100101; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b11101100; c = 8'b01000111; // Expected: {'sum': 193, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b11101100; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b11101010; c = 8'b01110001; // Expected: {'sum': 95, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b11101010; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b00001010; c = 8'b10010011; // Expected: {'sum': 71, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b00001010; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b01001011; c = 8'b10011011; // Expected: {'sum': 116, 'carry': 139}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b01001011; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01001110; c = 8'b11111111; // Expected: {'sum': 194, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01001110; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b11100010; c = 8'b00100010; // Expected: {'sum': 175, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b11100010; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01001001; c = 8'b00000110; // Expected: {'sum': 12, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01001001; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11111010; c = 8'b01101011; // Expected: {'sum': 135, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11111010; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b01101000; c = 8'b11111001; // Expected: {'sum': 239, 'carry': 120}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b01101000; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100111; b = 8'b11101001; c = 8'b11011101; // Expected: {'sum': 211, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100111; b = 8'b11101001; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b10001101; c = 8'b10011000; // Expected: {'sum': 108, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b10001101; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01101100; c = 8'b01110101; // Expected: {'sum': 118, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01101100; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b00000110; c = 8'b11110110; // Expected: {'sum': 44, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b00000110; c = 8'b11110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b01100011; c = 8'b11100000; // Expected: {'sum': 50, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b01100011; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b01101010; c = 8'b01111010; // Expected: {'sum': 99, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b01101010; c = 8'b01111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100100; b = 8'b10101000; c = 8'b11100100; // Expected: {'sum': 232, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100100; b = 8'b10101000; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b01000011; c = 8'b00001110; // Expected: {'sum': 245, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b01000011; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b11111001; c = 8'b01001110; // Expected: {'sum': 191, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b11111001; c = 8'b01001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100000; b = 8'b11101011; c = 8'b00000011; // Expected: {'sum': 8, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100000; b = 8'b11101011; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000100; b = 8'b00010100; c = 8'b11101001; // Expected: {'sum': 185, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000100; b = 8'b00010100; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b11000110; c = 8'b11001010; // Expected: {'sum': 39, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b11000110; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111100; b = 8'b11100011; c = 8'b10100100; // Expected: {'sum': 123, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111100; b = 8'b11100011; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01111011; c = 8'b00110100; // Expected: {'sum': 98, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01111011; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000100; b = 8'b10100010; c = 8'b00100101; // Expected: {'sum': 3, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000100; b = 8'b10100010; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b01101101; c = 8'b11011011; // Expected: {'sum': 47, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b01101101; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10111010; c = 8'b11011110; // Expected: {'sum': 119, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10111010; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 119, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00000111; c = 8'b01001111; // Expected: {'sum': 227, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00000111; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01111101; c = 8'b11011111; // Expected: {'sum': 156, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01111101; c = 8'b11011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10110100; c = 8'b10101110; // Expected: {'sum': 181, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10110100; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b11101001; c = 8'b00111000; // Expected: {'sum': 16, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b11101001; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b11010100; c = 8'b00100010; // Expected: {'sum': 237, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b11010100; c = 8'b00100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10000100; c = 8'b10110011; // Expected: {'sum': 214, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10000100; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 214, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00111011; c = 8'b11100101; // Expected: {'sum': 123, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00111011; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b11110001; c = 8'b01110010; // Expected: {'sum': 224, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b11110001; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b10110110; c = 8'b11000110; // Expected: {'sum': 247, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b10110110; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b10100011; c = 8'b11110010; // Expected: {'sum': 152, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b10100011; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b01110111; c = 8'b10011111; // Expected: {'sum': 9, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b01110111; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101110; b = 8'b10010110; c = 8'b01011110; // Expected: {'sum': 230, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101110; b = 8'b10010110; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b10000011; c = 8'b00001010; // Expected: {'sum': 125, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b10000011; c = 8'b00001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 125, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b01111110; c = 8'b00010001; // Expected: {'sum': 38, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b01111110; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b01110001; c = 8'b00001101; // Expected: {'sum': 60, 'carry': 65}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b01110001; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11010011; c = 8'b11111001; // Expected: {'sum': 38, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11010011; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 38, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b00011100; c = 8'b10101111; // Expected: {'sum': 93, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b00011100; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b00111000; c = 8'b00101100; // Expected: {'sum': 65, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b00111000; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b00010100; c = 8'b01010010; // Expected: {'sum': 98, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b00010100; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101010; b = 8'b00101011; c = 8'b11011100; // Expected: {'sum': 157, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101010; b = 8'b00101011; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 157, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b00010101; c = 8'b00100101; // Expected: {'sum': 137, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b00010101; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01111111; c = 8'b00101000; // Expected: {'sum': 209, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01111111; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b10011010; c = 8'b01001100; // Expected: {'sum': 228, 'carry': 26}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b10011010; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00110101; c = 8'b01100100; // Expected: {'sum': 61, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00110101; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11010000; c = 8'b00100011; // Expected: {'sum': 138, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11010000; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00001010; c = 8'b10111111; // Expected: {'sum': 209, 'carry': 46}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00001010; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b01001100; c = 8'b01011001; // Expected: {'sum': 118, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b01001100; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b00001001; c = 8'b00111101; // Expected: {'sum': 95, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b00001001; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b11001111; c = 8'b00111011; // Expected: {'sum': 222, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b11001111; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100011; b = 8'b11111011; c = 8'b11100011; // Expected: {'sum': 59, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100011; b = 8'b11111011; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b10111001; c = 8'b01001000; // Expected: {'sum': 83, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b10111001; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000000; b = 8'b11111100; c = 8'b11011100; // Expected: {'sum': 224, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000000; b = 8'b11111100; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 224, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b11111011; c = 8'b10000010; // Expected: {'sum': 191, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b11111011; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00001011; c = 8'b00000111; // Expected: {'sum': 65, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00001011; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10001000; c = 8'b11111001; // Expected: {'sum': 158, 'carry': 233}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10001000; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110001; b = 8'b10101110; c = 8'b10000100; // Expected: {'sum': 219, 'carry': 164}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110001; b = 8'b10101110; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 219, 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010011; b = 8'b11101111; c = 8'b10111111; // Expected: {'sum': 131, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010011; b = 8'b11101111; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01100101; c = 8'b01101101; // Expected: {'sum': 0, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01100101; c = 8'b01101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b10110011; c = 8'b10101001; // Expected: {'sum': 64, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b10110011; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10100001; c = 8'b10011011; // Expected: {'sum': 132, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10100001; c = 8'b10011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 132, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b10111100; c = 8'b11001111; // Expected: {'sum': 209, 'carry': 174}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b10111100; c = 8'b11001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111111; b = 8'b00010001; c = 8'b00001101; // Expected: {'sum': 227, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111111; b = 8'b00010001; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01001100; c = 8'b10011000; // Expected: {'sum': 58, 'carry': 204}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01001100; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 58, 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11101000; c = 8'b10110011; // Expected: {'sum': 19, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11101000; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b11110111; c = 8'b10010101; // Expected: {'sum': 14, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b11110111; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b01111101; c = 8'b00011110; // Expected: {'sum': 5, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b01111101; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111111; b = 8'b01101001; c = 8'b10101111; // Expected: {'sum': 185, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111111; b = 8'b01101001; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b10001101; c = 8'b01100100; // Expected: {'sum': 241, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b10001101; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b00101001; c = 8'b10000000; // Expected: {'sum': 77, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b00101001; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101011; b = 8'b00100001; c = 8'b10110111; // Expected: {'sum': 189, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101011; b = 8'b00100001; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b11001111; c = 8'b01010100; // Expected: {'sum': 175, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b11001111; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011010; b = 8'b10101110; c = 8'b01110010; // Expected: {'sum': 198, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011010; b = 8'b10101110; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 198, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b00101001; c = 8'b01001000; // Expected: {'sum': 76, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b00101001; c = 8'b01001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b00001011; c = 8'b00011001; // Expected: {'sum': 12, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b00001011; c = 8'b00011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b00110100; c = 8'b00111110; // Expected: {'sum': 18, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b00110100; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b01110101; c = 8'b01101011; // Expected: {'sum': 134, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b01110101; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00010011; c = 8'b11010001; // Expected: {'sum': 197, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00010011; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 197, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10101000; c = 8'b11010111; // Expected: {'sum': 53, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10101000; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01001010; c = 8'b10111101; // Expected: {'sum': 163, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01001010; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10100100; c = 8'b01101011; // Expected: {'sum': 71, 'carry': 168}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10100100; c = 8'b01101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 71, 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b01010100; c = 8'b11110111; // Expected: {'sum': 113, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b01010100; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001011; b = 8'b00111001; c = 8'b10100011; // Expected: {'sum': 145, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001011; b = 8'b00111001; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01100100; c = 8'b10001011; // Expected: {'sum': 239, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01100100; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b11101101; c = 8'b11101000; // Expected: {'sum': 120, 'carry': 237}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b11101101; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b10011111; c = 8'b11010101; // Expected: {'sum': 84, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b10011111; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11010011; c = 8'b11011101; // Expected: {'sum': 220, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11010011; c = 8'b11011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110000; b = 8'b11010100; c = 8'b00011111; // Expected: {'sum': 59, 'carry': 212}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110000; b = 8'b11010100; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b11111010; c = 8'b01000100; // Expected: {'sum': 178, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b11111010; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b00000001; c = 8'b01101001; // Expected: {'sum': 164, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b00000001; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b01010010; c = 8'b01100001; // Expected: {'sum': 116, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b01010010; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b10101101; c = 8'b10011100; // Expected: {'sum': 128, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b10101101; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b01110001; c = 8'b00000100; // Expected: {'sum': 225, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b01110001; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00100001; c = 8'b10100010; // Expected: {'sum': 138, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00100001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b11010001; c = 8'b00110000; // Expected: {'sum': 235, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b11010001; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 235, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b10000101; c = 8'b01010011; // Expected: {'sum': 36, 'carry': 211}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b10000101; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 36, 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10111111; c = 8'b11100011; // Expected: {'sum': 103, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10111111; c = 8'b11100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001100; b = 8'b10100000; c = 8'b00111110; // Expected: {'sum': 146, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001100; b = 8'b10100000; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 146, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b01100111; c = 8'b00101010; // Expected: {'sum': 77, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b01100111; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b11110001; c = 8'b10110110; // Expected: {'sum': 99, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b11110001; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b11000101; c = 8'b11101111; // Expected: {'sum': 28, 'carry': 231}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b11000101; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b01011011; c = 8'b00101010; // Expected: {'sum': 253, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b01011011; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b10110110; c = 8'b11000110; // Expected: {'sum': 140, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b10110110; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01010111; c = 8'b11111111; // Expected: {'sum': 64, 'carry': 255}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01010111; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b10110101; c = 8'b11110001; // Expected: {'sum': 40, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b10110101; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10000111; c = 8'b11110011; // Expected: {'sum': 79, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10000111; c = 8'b11110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10100110; c = 8'b00000111; // Expected: {'sum': 151, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10100110; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11100011; c = 8'b11100101; // Expected: {'sum': 100, 'carry': 227}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11100011; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b01111010; c = 8'b11000110; // Expected: {'sum': 89, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b01111010; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b11110000; c = 8'b01110000; // Expected: {'sum': 92, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b11110000; c = 8'b01110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11000101; c = 8'b11110010; // Expected: {'sum': 203, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11000101; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b10011001; c = 8'b10010000; // Expected: {'sum': 121, 'carry': 144}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b10011001; c = 8'b10010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b11111100; c = 8'b00110000; // Expected: {'sum': 52, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b11111100; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b00011000; c = 8'b01100010; // Expected: {'sum': 168, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b00011000; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b01001001; c = 8'b11011001; // Expected: {'sum': 159, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b01001001; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 159, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100010; b = 8'b11011101; c = 8'b10001111; // Expected: {'sum': 48, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100010; b = 8'b11011101; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 48, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00111000; c = 8'b11111110; // Expected: {'sum': 156, 'carry': 122}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00111000; c = 8'b11111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 156, 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011010; b = 8'b00011010; c = 8'b11000110; // Expected: {'sum': 70, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011010; b = 8'b00011010; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11101011; c = 8'b00000111; // Expected: {'sum': 223, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11101011; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 223, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011110; b = 8'b10100101; c = 8'b11010110; // Expected: {'sum': 45, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011110; b = 8'b10100101; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 45, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10001111; c = 8'b10001110; // Expected: {'sum': 23, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10001111; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b00100000; c = 8'b00011111; // Expected: {'sum': 221, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b00100000; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 221, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00001101; c = 8'b01100100; // Expected: {'sum': 37, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00001101; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 37, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101001; b = 8'b01001001; c = 8'b01001100; // Expected: {'sum': 108, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101001; b = 8'b01001001; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b10001001; c = 8'b10001100; // Expected: {'sum': 72, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b10001001; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b11101101; c = 8'b10110000; // Expected: {'sum': 75, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b11101101; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b01111111; c = 8'b01111111; // Expected: {'sum': 95, 'carry': 127}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b01111111; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00100010; c = 8'b01110110; // Expected: {'sum': 116, 'carry': 34}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00100010; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100110; b = 8'b10001100; c = 8'b00001011; // Expected: {'sum': 97, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100110; b = 8'b10001100; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000010; b = 8'b01101011; c = 8'b10001001; // Expected: {'sum': 160, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000010; b = 8'b01101011; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b11100110; c = 8'b11000001; // Expected: {'sum': 250, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b11100110; c = 8'b11000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b11101011; c = 8'b10000010; // Expected: {'sum': 21, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b11101011; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b01101010; c = 8'b01111100; // Expected: {'sum': 28, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b01101010; c = 8'b01111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111101; b = 8'b10110110; c = 8'b11001010; // Expected: {'sum': 1, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111101; b = 8'b10110110; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100111; b = 8'b00101001; c = 8'b01011110; // Expected: {'sum': 16, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100111; b = 8'b00101001; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 16, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00111111; c = 8'b10101011; // Expected: {'sum': 52, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00111111; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011001; b = 8'b11010110; c = 8'b11101011; // Expected: {'sum': 100, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011001; b = 8'b11010110; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b10011010; c = 8'b01011001; // Expected: {'sum': 178, 'carry': 89}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b10011010; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110000; b = 8'b11100101; c = 8'b11011000; // Expected: {'sum': 13, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110000; b = 8'b11100101; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b01111000; c = 8'b10011110; // Expected: {'sum': 216, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b01111000; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00011000; c = 8'b11010110; // Expected: {'sum': 61, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00011000; c = 8'b11010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10111011; c = 8'b01011111; // Expected: {'sum': 46, 'carry': 219}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10111011; c = 8'b01011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10110111; c = 8'b10001010; // Expected: {'sum': 169, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10110111; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01000010; c = 8'b11110001; // Expected: {'sum': 128, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01000010; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01110110; c = 8'b10101011; // Expected: {'sum': 240, 'carry': 47}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01110110; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b00011111; c = 8'b11110000; // Expected: {'sum': 90, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b00011111; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100101; b = 8'b01111010; c = 8'b00100100; // Expected: {'sum': 59, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100101; b = 8'b01111010; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b11101111; c = 8'b00011101; // Expected: {'sum': 203, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b11101111; c = 8'b00011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b00011101; c = 8'b10101110; // Expected: {'sum': 8, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b00011101; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b10011111; c = 8'b01010100; // Expected: {'sum': 189, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b10011111; c = 8'b01010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 189, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b11000110; c = 8'b01101001; // Expected: {'sum': 180, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b11000110; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b01111100; c = 8'b10101001; // Expected: {'sum': 118, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b01111100; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 118, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110100; b = 8'b11001111; c = 8'b01100100; // Expected: {'sum': 31, 'carry': 228}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110100; b = 8'b11001111; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00011101; c = 8'b01101100; // Expected: {'sum': 199, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00011101; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 199, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100101; b = 8'b00100110; c = 8'b00001001; // Expected: {'sum': 202, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100101; b = 8'b00100110; c = 8'b00001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b01011010; c = 8'b00101001; // Expected: {'sum': 52, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b01011010; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 52, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b00010110; c = 8'b10000011; // Expected: {'sum': 62, 'carry': 131}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b00010110; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b10001001; c = 8'b01100101; // Expected: {'sum': 114, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b10001001; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111110; b = 8'b10100001; c = 8'b00011110; // Expected: {'sum': 129, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111110; b = 8'b10100001; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b01011010; c = 8'b10011001; // Expected: {'sum': 110, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b01011010; c = 8'b10011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00001011; c = 8'b11011010; // Expected: {'sum': 150, 'carry': 75}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00001011; c = 8'b11011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110101; b = 8'b11011001; c = 8'b10001111; // Expected: {'sum': 35, 'carry': 221}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110101; b = 8'b11011001; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00001010; c = 8'b01111001; // Expected: {'sum': 128, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00001010; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10000001; c = 8'b10100110; // Expected: {'sum': 109, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10000001; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10001110; c = 8'b10001010; // Expected: {'sum': 3, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10001110; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01111011; c = 8'b00000100; // Expected: {'sum': 236, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01111011; c = 8'b00000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 236, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001100; b = 8'b01011000; c = 8'b11010101; // Expected: {'sum': 1, 'carry': 220}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001100; b = 8'b01011000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01001111; c = 8'b00100001; // Expected: {'sum': 84, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01001111; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b00100101; c = 8'b11100100; // Expected: {'sum': 151, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b00100101; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b11110000; c = 8'b01000100; // Expected: {'sum': 163, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b11110000; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b01101101; c = 8'b01111110; // Expected: {'sum': 163, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b01101101; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b11010001; c = 8'b11000011; // Expected: {'sum': 251, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b11010001; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 251, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b10010101; c = 8'b01011001; // Expected: {'sum': 6, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b10010101; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11011111; c = 8'b01001011; // Expected: {'sum': 249, 'carry': 79}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11011111; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b01111110; c = 8'b10111101; // Expected: {'sum': 94, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b01111110; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110110; b = 8'b01101100; c = 8'b00010111; // Expected: {'sum': 141, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110110; b = 8'b01101100; c = 8'b00010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010110; b = 8'b11010011; c = 8'b01111110; // Expected: {'sum': 123, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010110; b = 8'b11010011; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b00101100; c = 8'b00010101; // Expected: {'sum': 131, 'carry': 60}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b00101100; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b01100011; c = 8'b00100111; // Expected: {'sum': 172, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b01100011; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10000101; c = 8'b11011011; // Expected: {'sum': 247, 'carry': 137}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10000101; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b00011111; c = 8'b11000010; // Expected: {'sum': 73, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b00011111; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011111; b = 8'b00101010; c = 8'b00010001; // Expected: {'sum': 164, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011111; b = 8'b00101010; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11111000; c = 8'b00110111; // Expected: {'sum': 100, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11111000; c = 8'b00110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 100, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b00010100; c = 8'b11100010; // Expected: {'sum': 204, 'carry': 50}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b00010100; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00011011; c = 8'b10111101; // Expected: {'sum': 209, 'carry': 63}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00011011; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 209, 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b00000000; c = 8'b01111110; // Expected: {'sum': 106, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b00000000; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 106, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01000100; c = 8'b11101111; // Expected: {'sum': 211, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01000100; c = 8'b11101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 211, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000110; b = 8'b10001000; c = 8'b00101110; // Expected: {'sum': 96, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000110; b = 8'b10001000; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10011010; c = 8'b00011111; // Expected: {'sum': 8, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10011010; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01011011; c = 8'b00111100; // Expected: {'sum': 11, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01011011; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b01110001; c = 8'b01110110; // Expected: {'sum': 26, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b01110001; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 26, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b01000010; c = 8'b00101110; // Expected: {'sum': 2, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b01000010; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10110100; c = 8'b01100110; // Expected: {'sum': 9, 'carry': 246}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10110100; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b11000111; c = 8'b01100000; // Expected: {'sum': 79, 'carry': 224}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b11000111; c = 8'b01100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 79, 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111101; b = 8'b00110111; c = 8'b00100000; // Expected: {'sum': 42, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111101; b = 8'b00110111; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100110; b = 8'b00110001; c = 8'b01100110; // Expected: {'sum': 49, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100110; b = 8'b00110001; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b00001000; c = 8'b10110110; // Expected: {'sum': 201, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b00001000; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b11011110; c = 8'b00001111; // Expected: {'sum': 168, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b11011110; c = 8'b00001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011110; b = 8'b00000101; c = 8'b01111101; // Expected: {'sum': 230, 'carry': 29}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011110; b = 8'b00000101; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 230, 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b00111011; c = 8'b00001000; // Expected: {'sum': 123, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b00111011; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10101000; c = 8'b10110111; // Expected: {'sum': 139, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10101000; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 139, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b11111110; c = 8'b01011010; // Expected: {'sum': 6, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b11111110; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b01111011; c = 8'b11111000; // Expected: {'sum': 2, 'carry': 249}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b01111011; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b11111011; c = 8'b10010110; // Expected: {'sum': 228, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b11111011; c = 8'b10010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b10110010; c = 8'b00100100; // Expected: {'sum': 192, 'carry': 54}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b10110010; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010111; b = 8'b00000100; c = 8'b00111011; // Expected: {'sum': 232, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010111; b = 8'b00000100; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00111010; c = 8'b11100001; // Expected: {'sum': 150, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00111010; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 150, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b00100010; c = 8'b00010101; // Expected: {'sum': 136, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b00100010; c = 8'b00010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 136, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b01100001; c = 8'b01110110; // Expected: {'sum': 145, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b01100001; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011000; b = 8'b00100001; c = 8'b10001001; // Expected: {'sum': 240, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011000; b = 8'b00100001; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01100000; c = 8'b00100100; // Expected: {'sum': 17, 'carry': 100}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01100000; c = 8'b00100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110111; b = 8'b11111101; c = 8'b01110101; // Expected: {'sum': 255, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110111; b = 8'b11111101; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00010101; c = 8'b10000000; // Expected: {'sum': 207, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00010101; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b00111110; c = 8'b00011011; // Expected: {'sum': 180, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b00111110; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111111; b = 8'b10110110; c = 8'b00111110; // Expected: {'sum': 55, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111111; b = 8'b10110110; c = 8'b00111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001010; b = 8'b10111110; c = 8'b01111000; // Expected: {'sum': 204, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001010; b = 8'b10111110; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 204, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b10110110; c = 8'b01110100; // Expected: {'sum': 98, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b10110110; c = 8'b01110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110100; b = 8'b00111001; c = 8'b00011111; // Expected: {'sum': 210, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110100; b = 8'b00111001; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00010111; c = 8'b00001101; // Expected: {'sum': 75, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00010111; c = 8'b00001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 75, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01110010; c = 8'b11010111; // Expected: {'sum': 129, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01110010; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 129, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11010101; c = 8'b01010000; // Expected: {'sum': 160, 'carry': 85}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11010101; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 160, 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b01100011; c = 8'b11110000; // Expected: {'sum': 222, 'carry': 97}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b01100011; c = 8'b11110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 222, 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b00011010; c = 8'b10011100; // Expected: {'sum': 232, 'carry': 30}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b00011010; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b00000010; c = 8'b11111100; // Expected: {'sum': 77, 'carry': 178}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b00000010; c = 8'b11111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b01010100; c = 8'b01001100; // Expected: {'sum': 14, 'carry': 84}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b01010100; c = 8'b01001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01111101; c = 8'b11001110; // Expected: {'sum': 203, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01111101; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b10001001; c = 8'b00101000; // Expected: {'sum': 148, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b10001001; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 148, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11010001; c = 8'b11101100; // Expected: {'sum': 188, 'carry': 193}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11010001; c = 8'b11101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 188, 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111000; b = 8'b00110011; c = 8'b11101010; // Expected: {'sum': 33, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111000; b = 8'b00110011; c = 8'b11101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b01100010; c = 8'b00100001; // Expected: {'sum': 0, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b01100010; c = 8'b00100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b10011001; c = 8'b10100100; // Expected: {'sum': 96, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b10011001; c = 8'b10100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 96, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b10111110; c = 8'b11001011; // Expected: {'sum': 167, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b10111110; c = 8'b11001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b00100111; c = 8'b01111001; // Expected: {'sum': 74, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b00100111; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b11111010; c = 8'b00011011; // Expected: {'sum': 164, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b11111010; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b11000100; c = 8'b00110001; // Expected: {'sum': 9, 'carry': 244}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b11000100; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00011000; c = 8'b10001110; // Expected: {'sum': 30, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00011000; c = 8'b10001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b00101000; c = 8'b01100001; // Expected: {'sum': 164, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b00101000; c = 8'b01100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b10100010; c = 8'b00010010; // Expected: {'sum': 248, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b10100010; c = 8'b00010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100011; b = 8'b10000000; c = 8'b10000001; // Expected: {'sum': 162, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100011; b = 8'b10000000; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 162, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b01100110; c = 8'b10111010; // Expected: {'sum': 179, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b01100110; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111010; b = 8'b10011011; c = 8'b00101000; // Expected: {'sum': 9, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111010; b = 8'b10011011; c = 8'b00101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011011; b = 8'b00010110; c = 8'b00100111; // Expected: {'sum': 106, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011011; b = 8'b00010110; c = 8'b00100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 106, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10101001; c = 8'b11101011; // Expected: {'sum': 173, 'carry': 235}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10101001; c = 8'b11101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b10111010; c = 8'b00101001; // Expected: {'sum': 149, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b10111010; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 149, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111101; b = 8'b01000001; c = 8'b10111110; // Expected: {'sum': 66, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111101; b = 8'b01000001; c = 8'b10111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b01001111; c = 8'b11011110; // Expected: {'sum': 35, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b01001111; c = 8'b11011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b00010100; c = 8'b10100111; // Expected: {'sum': 68, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b00010100; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b00011101; c = 8'b10110101; // Expected: {'sum': 175, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b00011101; c = 8'b10110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100010; b = 8'b10110001; c = 8'b10011100; // Expected: {'sum': 207, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100010; b = 8'b10110001; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 207, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000110; b = 8'b11001000; c = 8'b00001000; // Expected: {'sum': 134, 'carry': 72}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000110; b = 8'b11001000; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110000; b = 8'b00100001; c = 8'b10001100; // Expected: {'sum': 29, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110000; b = 8'b00100001; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b10010101; c = 8'b11110010; // Expected: {'sum': 34, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b10010101; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 34, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000101; b = 8'b01010000; c = 8'b10010001; // Expected: {'sum': 68, 'carry': 145}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000101; b = 8'b01010000; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011100; b = 8'b10101001; c = 8'b00000010; // Expected: {'sum': 247, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011100; b = 8'b10101001; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b10000000; c = 8'b10110001; // Expected: {'sum': 17, 'carry': 160}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b10000000; c = 8'b10110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11101010; c = 8'b10001011; // Expected: {'sum': 84, 'carry': 171}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11101010; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 84, 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001001; b = 8'b00100010; c = 8'b11011001; // Expected: {'sum': 178, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001001; b = 8'b00100010; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 178, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100000; b = 8'b00111110; c = 8'b10011010; // Expected: {'sum': 4, 'carry': 186}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100000; b = 8'b00111110; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b10111010; c = 8'b10111000; // Expected: {'sum': 143, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b10111010; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 143, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b00001101; c = 8'b11110100; // Expected: {'sum': 145, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b00001101; c = 8'b11110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b10110000; c = 8'b00011110; // Expected: {'sum': 53, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b10110000; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11110111; c = 8'b10101100; // Expected: {'sum': 234, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11110111; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000111; b = 8'b10111000; c = 8'b01110001; // Expected: {'sum': 206, 'carry': 49}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000111; b = 8'b10111000; c = 8'b01110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 206, 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010000; b = 8'b10110111; c = 8'b01010110; // Expected: {'sum': 241, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010000; b = 8'b10110111; c = 8'b01010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10100100; c = 8'b10001101; // Expected: {'sum': 175, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10100100; c = 8'b10001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101000; b = 8'b11000101; c = 8'b00111100; // Expected: {'sum': 17, 'carry': 236}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101000; b = 8'b11000101; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b11010010; c = 8'b11111010; // Expected: {'sum': 121, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b11010010; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b00000011; c = 8'b00111101; // Expected: {'sum': 183, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b00000011; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110000; b = 8'b01000000; c = 8'b10010011; // Expected: {'sum': 163, 'carry': 80}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110000; b = 8'b01000000; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 163, 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b11011111; c = 8'b10101110; // Expected: {'sum': 120, 'carry': 143}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b11011111; c = 8'b10101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 120, 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01011100; c = 8'b01001010; // Expected: {'sum': 92, 'carry': 74}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01011100; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b01010001; c = 8'b00011010; // Expected: {'sum': 185, 'carry': 82}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b01010001; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10110111; c = 8'b00101111; // Expected: {'sum': 185, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10110111; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b10100111; c = 8'b00000111; // Expected: {'sum': 216, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b10100111; c = 8'b00000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 216, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b10000001; c = 8'b11001110; // Expected: {'sum': 15, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b10000001; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01011011; c = 8'b01111101; // Expected: {'sum': 131, 'carry': 125}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01011011; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 131, 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011111; b = 8'b10001111; c = 8'b01110011; // Expected: {'sum': 35, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011111; b = 8'b10001111; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01001111; c = 8'b01000100; // Expected: {'sum': 201, 'carry': 70}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01001111; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001110; b = 8'b10010100; c = 8'b00110101; // Expected: {'sum': 47, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001110; b = 8'b10010100; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 47, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b01100101; c = 8'b01111111; // Expected: {'sum': 151, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b01100101; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 151, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111001; b = 8'b11011110; c = 8'b00111101; // Expected: {'sum': 90, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111001; b = 8'b11011110; c = 8'b00111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b01010110; c = 8'b11101000; // Expected: {'sum': 55, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b01010110; c = 8'b11101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010001; b = 8'b10101111; c = 8'b00100110; // Expected: {'sum': 152, 'carry': 39}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010001; b = 8'b10101111; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01101110; c = 8'b01001010; // Expected: {'sum': 140, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01101110; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00100110; c = 8'b01111000; // Expected: {'sum': 172, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00100110; c = 8'b01111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 172, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b01101111; c = 8'b11011000; // Expected: {'sum': 33, 'carry': 222}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b01101111; c = 8'b11011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100010; b = 8'b00010100; c = 8'b11001001; // Expected: {'sum': 127, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100010; b = 8'b00010100; c = 8'b11001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000101; b = 8'b00001001; c = 8'b11000110; // Expected: {'sum': 10, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000101; b = 8'b00001001; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b11101110; c = 8'b00110011; // Expected: {'sum': 181, 'carry': 106}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b11101110; c = 8'b00110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 181, 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b01100100; c = 8'b10010111; // Expected: {'sum': 103, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b01100100; c = 8'b10010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000100; b = 8'b01110101; c = 8'b10001111; // Expected: {'sum': 62, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000100; b = 8'b01110101; c = 8'b10001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b10110110; c = 8'b11111111; // Expected: {'sum': 245, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b10110110; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011100; b = 8'b01001011; c = 8'b01110101; // Expected: {'sum': 226, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011100; b = 8'b01001011; c = 8'b01110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111110; b = 8'b10000100; c = 8'b01011011; // Expected: {'sum': 161, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111110; b = 8'b10000100; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b10001101; c = 8'b11110001; // Expected: {'sum': 194, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b10001101; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b10010001; c = 8'b11100010; // Expected: {'sum': 86, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b10010001; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011000; b = 8'b01101000; c = 8'b10100111; // Expected: {'sum': 23, 'carry': 232}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011000; b = 8'b01101000; c = 8'b10100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 23, 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b00101111; c = 8'b01110010; // Expected: {'sum': 29, 'carry': 98}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b00101111; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b01010011; c = 8'b00011000; // Expected: {'sum': 140, 'carry': 83}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b01010011; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010000; b = 8'b00011000; c = 8'b10000000; // Expected: {'sum': 200, 'carry': 16}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010000; b = 8'b00011000; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b10110001; c = 8'b00001000; // Expected: {'sum': 167, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b10110001; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 167, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b01110110; c = 8'b10010100; // Expected: {'sum': 94, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b01110110; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11010011; c = 8'b10111111; // Expected: {'sum': 237, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11010011; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 237, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b10100000; c = 8'b10000110; // Expected: {'sum': 101, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b10100000; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b10000101; c = 8'b00001011; // Expected: {'sum': 57, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b10000101; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b11001111; c = 8'b00011110; // Expected: {'sum': 50, 'carry': 207}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b11001111; c = 8'b00011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 50, 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b01110111; c = 8'b11111001; // Expected: {'sum': 171, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b01110111; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000111; b = 8'b11010101; c = 8'b01100110; // Expected: {'sum': 116, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000111; b = 8'b11010101; c = 8'b01100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b01001010; c = 8'b00101101; // Expected: {'sum': 242, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b01001010; c = 8'b00101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b00010000; c = 8'b10000100; // Expected: {'sum': 93, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b00010000; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 93, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00001111; c = 8'b00000110; // Expected: {'sum': 41, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00001111; c = 8'b00000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11000110; c = 8'b01001111; // Expected: {'sum': 31, 'carry': 198}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11000110; c = 8'b01001111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 31, 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010011; b = 8'b01011001; c = 8'b01011011; // Expected: {'sum': 145, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010011; b = 8'b01011001; c = 8'b01011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 145, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b00100110; c = 8'b11100100; // Expected: {'sum': 141, 'carry': 102}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b00100110; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 141, 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101010; b = 8'b10111000; c = 8'b01011101; // Expected: {'sum': 15, 'carry': 248}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101010; b = 8'b10111000; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011000; b = 8'b11111001; c = 8'b11000000; // Expected: {'sum': 33, 'carry': 216}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011000; b = 8'b11111001; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 33, 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110100; b = 8'b00110100; c = 8'b10111111; // Expected: {'sum': 191, 'carry': 52}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110100; b = 8'b00110100; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10110100; c = 8'b10110011; // Expected: {'sum': 8, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10110100; c = 8'b10110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b10000111; c = 8'b00101011; // Expected: {'sum': 194, 'carry': 47}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b10000111; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100110; b = 8'b00100101; c = 8'b01111001; // Expected: {'sum': 122, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100110; b = 8'b00100101; c = 8'b01111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 122, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b10010011; c = 8'b11000100; // Expected: {'sum': 173, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b10010011; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b00001011; c = 8'b01100100; // Expected: {'sum': 140, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b00001011; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000111; b = 8'b00001111; c = 8'b10000010; // Expected: {'sum': 202, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000111; b = 8'b00001111; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110010; b = 8'b00010111; c = 8'b00010001; // Expected: {'sum': 180, 'carry': 19}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110010; b = 8'b00010111; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10000000; c = 8'b00000001; // Expected: {'sum': 110, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10000000; c = 8'b00000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 110, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100101; b = 8'b11011100; c = 8'b11010001; // Expected: {'sum': 40, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100101; b = 8'b11011100; c = 8'b11010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001111; b = 8'b10110010; c = 8'b11100010; // Expected: {'sum': 95, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001111; b = 8'b10110010; c = 8'b11100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00011010; c = 8'b01100101; // Expected: {'sum': 114, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00011010; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 114, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b11001101; c = 8'b01011001; // Expected: {'sum': 86, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b11001101; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 86, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b10111110; c = 8'b01001011; // Expected: {'sum': 185, 'carry': 78}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b10111110; c = 8'b01001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110110; b = 8'b00000110; c = 8'b10011100; // Expected: {'sum': 44, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110110; b = 8'b00000110; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 44, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b11111010; c = 8'b01011110; // Expected: {'sum': 69, 'carry': 250}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b11111010; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 69, 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b11010110; c = 8'b10101100; // Expected: {'sum': 177, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b11010110; c = 8'b10101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b00110101; c = 8'b00011010; // Expected: {'sum': 126, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b00110101; c = 8'b00011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101111; b = 8'b00000101; c = 8'b01011100; // Expected: {'sum': 54, 'carry': 77}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101111; b = 8'b00000101; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b11010111; c = 8'b01100111; // Expected: {'sum': 1, 'carry': 247}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b11010111; c = 8'b01100111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010111; b = 8'b11011110; c = 8'b00111000; // Expected: {'sum': 177, 'carry': 94}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010111; b = 8'b11011110; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 177, 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b00001101; c = 8'b01000001; // Expected: {'sum': 95, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b00001101; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010101; b = 8'b01110111; c = 8'b11010111; // Expected: {'sum': 245, 'carry': 87}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010101; b = 8'b01110111; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010101; b = 8'b11111010; c = 8'b10000110; // Expected: {'sum': 233, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010101; b = 8'b11111010; c = 8'b10000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b00111101; c = 8'b10111011; // Expected: {'sum': 254, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b00111101; c = 8'b10111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 254, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011111; b = 8'b10001101; c = 8'b10110000; // Expected: {'sum': 98, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011111; b = 8'b10001101; c = 8'b10110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101011; b = 8'b00111010; c = 8'b11100100; // Expected: {'sum': 53, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101011; b = 8'b00111010; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b01001101; c = 8'b11110010; // Expected: {'sum': 137, 'carry': 118}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b01001101; c = 8'b11110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110101; b = 8'b11010111; c = 8'b00100110; // Expected: {'sum': 196, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110101; b = 8'b11010111; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 196, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b01100001; c = 8'b00110101; // Expected: {'sum': 0, 'carry': 117}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b01100001; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b11011110; c = 8'b01001101; // Expected: {'sum': 40, 'carry': 223}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b11011110; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001101; b = 8'b00001001; c = 8'b00111011; // Expected: {'sum': 127, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001101; b = 8'b00001001; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 127, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b10011001; c = 8'b10111111; // Expected: {'sum': 108, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b10011001; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 108, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010010; b = 8'b01101011; c = 8'b10001001; // Expected: {'sum': 240, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010010; b = 8'b01101011; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 240, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101100; b = 8'b10010001; c = 8'b01111111; // Expected: {'sum': 2, 'carry': 253}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101100; b = 8'b10010001; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110010; b = 8'b11100010; c = 8'b10000101; // Expected: {'sum': 21, 'carry': 226}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110010; b = 8'b11100010; c = 8'b10000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010011; b = 8'b10011001; c = 8'b11001100; // Expected: {'sum': 70, 'carry': 153}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010011; b = 8'b10011001; c = 8'b11001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 70, 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b10111001; c = 8'b10110110; // Expected: {'sum': 248, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b10111001; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 248, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01001100; c = 8'b01011101; // Expected: {'sum': 105, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01001100; c = 8'b01011101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b10011000; c = 8'b01101001; // Expected: {'sum': 213, 'carry': 40}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b10011000; c = 8'b01101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b10001000; c = 8'b10101000; // Expected: {'sum': 99, 'carry': 136}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b10001000; c = 8'b10101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110011; b = 8'b10101000; c = 8'b00001110; // Expected: {'sum': 213, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110011; b = 8'b10101000; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010100; b = 8'b00001010; c = 8'b10001010; // Expected: {'sum': 212, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010100; b = 8'b00001010; c = 8'b10001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110101; b = 8'b01101011; c = 8'b01010000; // Expected: {'sum': 142, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110101; b = 8'b01101011; c = 8'b01010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101010; b = 8'b11100100; c = 8'b00000010; // Expected: {'sum': 76, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101010; b = 8'b11100100; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110110; b = 8'b11011110; c = 8'b01000001; // Expected: {'sum': 233, 'carry': 86}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110110; b = 8'b11011110; c = 8'b01000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 233, 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00110101; c = 8'b01010111; // Expected: {'sum': 234, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00110101; c = 8'b01010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110111; b = 8'b01100001; c = 8'b10101101; // Expected: {'sum': 123, 'carry': 165}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110111; b = 8'b01100001; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 123, 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b00011100; c = 8'b00011000; // Expected: {'sum': 76, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b00011100; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 76, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011011; b = 8'b11100111; c = 8'b10010011; // Expected: {'sum': 239, 'carry': 147}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011011; b = 8'b11100111; c = 8'b10010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00010111; c = 8'b10011100; // Expected: {'sum': 137, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00010111; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 137, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b01001101; c = 8'b10110110; // Expected: {'sum': 49, 'carry': 206}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b01001101; c = 8'b10110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 49, 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10110100; c = 8'b00001110; // Expected: {'sum': 175, 'carry': 20}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10110100; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 175, 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b10101111; c = 8'b01100010; // Expected: {'sum': 212, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b10101111; c = 8'b01100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100001; b = 8'b00111010; c = 8'b11100101; // Expected: {'sum': 126, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100001; b = 8'b00111010; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00111010; c = 8'b10101111; // Expected: {'sum': 180, 'carry': 43}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00111010; c = 8'b10101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 180, 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101011; b = 8'b01101011; c = 8'b10111000; // Expected: {'sum': 184, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101011; b = 8'b01101011; c = 8'b10111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001101; b = 8'b00010010; c = 8'b01010010; // Expected: {'sum': 205, 'carry': 18}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001101; b = 8'b00010010; c = 8'b01010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111000; b = 8'b01011100; c = 8'b11100101; // Expected: {'sum': 193, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111000; b = 8'b01011100; c = 8'b11100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b10011101; c = 8'b00101100; // Expected: {'sum': 217, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b10011101; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 217, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b01100011; c = 8'b11010101; // Expected: {'sum': 19, 'carry': 229}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b01100011; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000111; b = 8'b10000011; c = 8'b00000101; // Expected: {'sum': 1, 'carry': 135}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000111; b = 8'b10000011; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b00111110; c = 8'b00101111; // Expected: {'sum': 82, 'carry': 47}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b00111110; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b11101001; c = 8'b10110111; // Expected: {'sum': 64, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b11101001; c = 8'b10110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000000; b = 8'b00110001; c = 8'b11011001; // Expected: {'sum': 232, 'carry': 17}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000000; b = 8'b00110001; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 232, 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b01100001; c = 8'b11011011; // Expected: {'sum': 128, 'carry': 123}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b01100001; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 128, 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11101011; c = 8'b00111011; // Expected: {'sum': 77, 'carry': 187}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11101011; c = 8'b00111011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b00100010; c = 8'b00100110; // Expected: {'sum': 171, 'carry': 38}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b00100010; c = 8'b00100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b01110100; c = 8'b00111100; // Expected: {'sum': 18, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b01110100; c = 8'b00111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b11111001; c = 8'b00000101; // Expected: {'sum': 68, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b11111001; c = 8'b00000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111100; b = 8'b00111110; c = 8'b01011100; // Expected: {'sum': 158, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111100; b = 8'b00111110; c = 8'b01011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b10110000; c = 8'b01000111; // Expected: {'sum': 92, 'carry': 163}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b10110000; c = 8'b01000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 92, 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010100; b = 8'b11111010; c = 8'b11100001; // Expected: {'sum': 15, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010100; b = 8'b11111010; c = 8'b11100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10011100; c = 8'b01101100; // Expected: {'sum': 105, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10011100; c = 8'b01101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 105, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010110; b = 8'b10000011; c = 8'b10001000; // Expected: {'sum': 29, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010110; b = 8'b10000011; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 29, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010110; b = 8'b01101011; c = 8'b01101110; // Expected: {'sum': 83, 'carry': 110}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010110; b = 8'b01101011; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 83, 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001111; b = 8'b11110001; c = 8'b11010111; // Expected: {'sum': 169, 'carry': 215}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001111; b = 8'b11110001; c = 8'b11010111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b00010001; c = 8'b11001110; // Expected: {'sum': 130, 'carry': 93}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b00010001; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b01011010; c = 8'b10111101; // Expected: {'sum': 53, 'carry': 218}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b01011010; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 53, 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000100; b = 8'b10001010; c = 8'b01000101; // Expected: {'sum': 203, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000100; b = 8'b10001010; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000110; b = 8'b10110110; c = 8'b00100101; // Expected: {'sum': 21, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000110; b = 8'b10110110; c = 8'b00100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 21, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110010; b = 8'b00101100; c = 8'b10111111; // Expected: {'sum': 161, 'carry': 62}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110010; b = 8'b00101100; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b01101000; c = 8'b11000011; // Expected: {'sum': 112, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b01101000; c = 8'b11000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b00110111; c = 8'b00010100; // Expected: {'sum': 234, 'carry': 21}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b00110111; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 234, 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01001010; c = 8'b10101011; // Expected: {'sum': 255, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01001010; c = 8'b10101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 255, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b01000010; c = 8'b11111010; // Expected: {'sum': 19, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b01000010; c = 8'b11111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101111; b = 8'b10100000; c = 8'b11000010; // Expected: {'sum': 205, 'carry': 162}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101111; b = 8'b10100000; c = 8'b11000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 205, 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111010; b = 8'b00110010; c = 8'b01000010; // Expected: {'sum': 138, 'carry': 114}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111010; b = 8'b00110010; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 138, 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011101; b = 8'b01111010; c = 8'b00111001; // Expected: {'sum': 30, 'carry': 121}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011101; b = 8'b01111010; c = 8'b00111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 30, 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11100101; c = 8'b10010010; // Expected: {'sum': 68, 'carry': 179}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11100101; c = 8'b10010010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 68, 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b01010111; c = 8'b11110111; // Expected: {'sum': 140, 'carry': 119}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b01010111; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100000; b = 8'b00011000; c = 8'b11011100; // Expected: {'sum': 228, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100000; b = 8'b00011000; c = 8'b11011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 228, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111100; b = 8'b10101101; c = 8'b00000010; // Expected: {'sum': 19, 'carry': 172}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111100; b = 8'b10101101; c = 8'b00000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 19, 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001110; b = 8'b11100010; c = 8'b00111000; // Expected: {'sum': 212, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001110; b = 8'b11100010; c = 8'b00111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 212, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101101; b = 8'b11000001; c = 8'b10010100; // Expected: {'sum': 56, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101101; b = 8'b11000001; c = 8'b10010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 56, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110111; b = 8'b11010110; c = 8'b10011110; // Expected: {'sum': 191, 'carry': 214}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110111; b = 8'b11010110; c = 8'b10011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 191, 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01011001; c = 8'b11001110; // Expected: {'sum': 63, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01011001; c = 8'b11001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b00000000; c = 8'b10011100; // Expected: {'sum': 28, 'carry': 128}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b00000000; c = 8'b10011100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b10111111; c = 8'b01110010; // Expected: {'sum': 99, 'carry': 190}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b10111111; c = 8'b01110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 99, 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001111; b = 8'b10000111; c = 8'b11110101; // Expected: {'sum': 61, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001111; b = 8'b10000111; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 61, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001000; b = 8'b01000100; c = 8'b10001100; // Expected: {'sum': 192, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001000; b = 8'b01000100; c = 8'b10001100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100011; b = 8'b10110101; c = 8'b00010110; // Expected: {'sum': 64, 'carry': 183}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100011; b = 8'b10110101; c = 8'b00010110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 64, 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01000000; c = 8'b00010001; // Expected: {'sum': 170, 'carry': 81}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01000000; c = 8'b00010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011011; b = 8'b00011111; c = 8'b10000011; // Expected: {'sum': 135, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011011; b = 8'b00011111; c = 8'b10000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 135, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001100; b = 8'b01111111; c = 8'b00101011; // Expected: {'sum': 152, 'carry': 111}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001100; b = 8'b01111111; c = 8'b00101011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 152, 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00000111; c = 8'b00110010; // Expected: {'sum': 192, 'carry': 55}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00000111; c = 8'b00110010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 192, 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000001; b = 8'b01110000; c = 8'b10000100; // Expected: {'sum': 245, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000001; b = 8'b01110000; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00101001; c = 8'b11111000; // Expected: {'sum': 77, 'carry': 184}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00101001; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 77, 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111100; b = 8'b00110001; c = 8'b01000010; // Expected: {'sum': 15, 'carry': 112}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111100; b = 8'b00110001; c = 8'b01000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10100000; c = 8'b10100011; // Expected: {'sum': 170, 'carry': 161}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10100000; c = 8'b10100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 170, 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101110; b = 8'b01101101; c = 8'b01100100; // Expected: {'sum': 103, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101110; b = 8'b01101101; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 103, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011110; b = 8'b01100110; c = 8'b00111010; // Expected: {'sum': 130, 'carry': 126}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011110; b = 8'b01100110; c = 8'b00111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 130, 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b10111001; c = 8'b01111111; // Expected: {'sum': 231, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b10111001; c = 8'b01111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101011; b = 8'b11101010; c = 8'b00001000; // Expected: {'sum': 73, 'carry': 170}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101011; b = 8'b11101010; c = 8'b00001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 73, 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000001; b = 8'b11110111; c = 8'b00110101; // Expected: {'sum': 67, 'carry': 181}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000001; b = 8'b11110111; c = 8'b00110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 67, 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111000; b = 8'b00101011; c = 8'b01011001; // Expected: {'sum': 202, 'carry': 57}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111000; b = 8'b00101011; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 202, 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b10111111; c = 8'b01101000; // Expected: {'sum': 126, 'carry': 169}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b10111111; c = 8'b01101000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 126, 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001101; b = 8'b00011111; c = 8'b11000000; // Expected: {'sum': 210, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001101; b = 8'b00011111; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 210, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101000; b = 8'b01100100; c = 8'b10011111; // Expected: {'sum': 147, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101000; b = 8'b01100100; c = 8'b10011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111001; b = 8'b10101001; c = 8'b01100101; // Expected: {'sum': 245, 'carry': 41}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111001; b = 8'b10101001; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 245, 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000010; b = 8'b01001111; c = 8'b11000111; // Expected: {'sum': 74, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000010; b = 8'b01001111; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 74, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010010; b = 8'b11101010; c = 8'b00101100; // Expected: {'sum': 20, 'carry': 234}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010010; b = 8'b11101010; c = 8'b00101100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001011; b = 8'b00010000; c = 8'b11001010; // Expected: {'sum': 17, 'carry': 202}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001011; b = 8'b00010000; c = 8'b11001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10100111; c = 8'b01011110; // Expected: {'sum': 113, 'carry': 142}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10100111; c = 8'b01011110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111111; b = 8'b11001111; c = 8'b01011001; // Expected: {'sum': 169, 'carry': 95}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111111; b = 8'b11001111; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 169, 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110011; b = 8'b10101111; c = 8'b01000110; // Expected: {'sum': 90, 'carry': 167}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110011; b = 8'b10101111; c = 8'b01000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 90, 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b10100110; c = 8'b11110001; // Expected: {'sum': 241, 'carry': 166}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b10100110; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011000; b = 8'b11100101; c = 8'b11011011; // Expected: {'sum': 166, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011000; b = 8'b11100101; c = 8'b11011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 166, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001001; b = 8'b10111101; c = 8'b11000101; // Expected: {'sum': 241, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001001; b = 8'b10111101; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 241, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010100; b = 8'b01001100; c = 8'b10100001; // Expected: {'sum': 57, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010100; b = 8'b01001100; c = 8'b10100001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 57, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111110; b = 8'b00101001; c = 8'b11110101; // Expected: {'sum': 98, 'carry': 189}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111110; b = 8'b00101001; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 98, 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10000000; b = 8'b10000110; c = 8'b00101111; // Expected: {'sum': 41, 'carry': 134}
        #10;
        $display("Test %0d: Inputs: a = 8'b10000000; b = 8'b10000110; c = 8'b00101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 41, 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111000; b = 8'b10100010; c = 8'b00100000; // Expected: {'sum': 186, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111000; b = 8'b10100010; c = 8'b00100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 186, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00100011; c = 8'b10100110; // Expected: {'sum': 140, 'carry': 35}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00100011; c = 8'b10100110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 140, 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b10011110; c = 8'b10111101; // Expected: {'sum': 171, 'carry': 156}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b10011110; c = 8'b10111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 171, 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101111; b = 8'b10101000; c = 8'b01101111; // Expected: {'sum': 40, 'carry': 239}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101111; b = 8'b10101000; c = 8'b01101111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b11000100; c = 8'b11000000; // Expected: {'sum': 55, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b11000100; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 55, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001000; b = 8'b11001011; c = 8'b10101001; // Expected: {'sum': 42, 'carry': 201}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001000; b = 8'b11001011; c = 8'b10101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 42, 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000001; b = 8'b01001010; c = 8'b11111111; // Expected: {'sum': 116, 'carry': 203}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000001; b = 8'b01001010; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 116, 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101010; b = 8'b01101101; c = 8'b00101010; // Expected: {'sum': 109, 'carry': 42}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101010; b = 8'b01101101; c = 8'b00101010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 109, 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00001001; b = 8'b00000011; c = 8'b00011011; // Expected: {'sum': 17, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 8'b00001001; b = 8'b00000011; c = 8'b00011011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 17, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111010; b = 8'b10101100; c = 8'b01100101; // Expected: {'sum': 243, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111010; b = 8'b10101100; c = 8'b01100101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 243, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100001; b = 8'b10111111; c = 8'b01010101; // Expected: {'sum': 11, 'carry': 245}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100001; b = 8'b10111111; c = 8'b01010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101001; b = 8'b11110010; c = 8'b10110100; // Expected: {'sum': 239, 'carry': 176}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101001; b = 8'b11110010; c = 8'b10110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 239, 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110110; b = 8'b10010100; c = 8'b10000001; // Expected: {'sum': 35, 'carry': 148}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110110; b = 8'b10010100; c = 8'b10000001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 35, 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001110; b = 8'b01111001; c = 8'b10001000; // Expected: {'sum': 63, 'carry': 200}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001110; b = 8'b01111001; c = 8'b10001000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 63, 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010110; b = 8'b11010011; c = 8'b10100010; // Expected: {'sum': 231, 'carry': 146}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010110; b = 8'b11010011; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 231, 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b10001010; c = 8'b10101101; // Expected: {'sum': 242, 'carry': 141}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b10001010; c = 8'b10101101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 242, 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011101; b = 8'b00110001; c = 8'b01101110; // Expected: {'sum': 66, 'carry': 61}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011101; b = 8'b00110001; c = 8'b01101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 66, 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010000; b = 8'b01010001; c = 8'b11100100; // Expected: {'sum': 101, 'carry': 208}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010000; b = 8'b01010001; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b11010110; c = 8'b01110011; // Expected: {'sum': 111, 'carry': 210}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b11010110; c = 8'b01110011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 111, 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b00110110; c = 8'b10111100; // Expected: {'sum': 121, 'carry': 182}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b00110110; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 121, 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b11001100; c = 8'b01011001; // Expected: {'sum': 185, 'carry': 76}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b11001100; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 185, 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01110001; b = 8'b00110001; c = 8'b01111110; // Expected: {'sum': 62, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b01110001; b = 8'b00110001; c = 8'b01111110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000000; b = 8'b11011100; c = 8'b01111101; // Expected: {'sum': 225, 'carry': 92}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000000; b = 8'b11011100; c = 8'b01111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 225, 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110101; b = 8'b00001000; c = 8'b11010101; // Expected: {'sum': 40, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110101; b = 8'b00001000; c = 8'b11010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011011; b = 8'b10111001; c = 8'b00000011; // Expected: {'sum': 97, 'carry': 155}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011011; b = 8'b10111001; c = 8'b00000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 97, 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001000; b = 8'b00001100; c = 8'b01000101; // Expected: {'sum': 193, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001000; b = 8'b00001100; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 193, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b00010101; c = 8'b10001001; // Expected: {'sum': 208, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b00010101; c = 8'b10001001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 208, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01011010; b = 8'b00000100; c = 8'b10001011; // Expected: {'sum': 213, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 8'b01011010; b = 8'b00000100; c = 8'b10001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 213, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100101; b = 8'b00000011; c = 8'b10011000; // Expected: {'sum': 62, 'carry': 129}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100101; b = 8'b00000011; c = 8'b10011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 62, 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11110000; c = 8'b01011000; // Expected: {'sum': 183, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11110000; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 183, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100011; b = 8'b10101101; c = 8'b00010100; // Expected: {'sum': 218, 'carry': 37}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100011; b = 8'b10101101; c = 8'b00010100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11010101; b = 8'b00010110; c = 8'b11000101; // Expected: {'sum': 6, 'carry': 213}
        #10;
        $display("Test %0d: Inputs: a = 8'b11010101; b = 8'b00010110; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011001; b = 8'b01100110; c = 8'b00001110; // Expected: {'sum': 113, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011001; b = 8'b01100110; c = 8'b00001110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 113, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010101; b = 8'b10010010; c = 8'b11000110; // Expected: {'sum': 65, 'carry': 150}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010101; b = 8'b10010010; c = 8'b11000110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 65, 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010111; b = 8'b10101110; c = 8'b10111111; // Expected: {'sum': 134, 'carry': 191}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010111; b = 8'b10101110; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 134, 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011111; b = 8'b11000000; c = 8'b01100100; // Expected: {'sum': 187, 'carry': 68}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011111; b = 8'b11000000; c = 8'b01100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 187, 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001010; b = 8'b01111100; c = 8'b11111101; // Expected: {'sum': 203, 'carry': 124}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001010; b = 8'b01111100; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 203, 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111011; b = 8'b01011011; c = 8'b10111100; // Expected: {'sum': 28, 'carry': 251}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111011; b = 8'b01011011; c = 8'b10111100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 28, 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001011; b = 8'b00010110; c = 8'b10010101; // Expected: {'sum': 200, 'carry': 23}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001011; b = 8'b00010110; c = 8'b10010101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11111110; b = 8'b00111100; c = 8'b11010000; // Expected: {'sum': 18, 'carry': 252}
        #10;
        $display("Test %0d: Inputs: a = 8'b11111110; b = 8'b00111100; c = 8'b11010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 18, 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00010111; c = 8'b00001011; // Expected: {'sum': 101, 'carry': 27}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00010111; c = 8'b00001011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 101, 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110011; b = 8'b01110001; c = 8'b00100011; // Expected: {'sum': 161, 'carry': 115}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110011; b = 8'b01110001; c = 8'b00100011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 161, 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10110001; b = 8'b00011000; c = 8'b01001010; // Expected: {'sum': 227, 'carry': 24}
        #10;
        $display("Test %0d: Inputs: a = 8'b10110001; b = 8'b00011000; c = 8'b01001010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010001; b = 8'b11111110; c = 8'b01011001; // Expected: {'sum': 54, 'carry': 217}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010001; b = 8'b11111110; c = 8'b01011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 54, 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001010; b = 8'b00101001; c = 8'b01001101; // Expected: {'sum': 174, 'carry': 73}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001010; b = 8'b00101001; c = 8'b01001101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 174, 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01001100; b = 8'b11111001; c = 8'b00010000; // Expected: {'sum': 165, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b01001100; b = 8'b11111001; c = 8'b00010000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101100; b = 8'b00000110; c = 8'b10000100; // Expected: {'sum': 46, 'carry': 132}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101100; b = 8'b00000110; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 46, 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10111011; b = 8'b01001100; c = 8'b01010011; // Expected: {'sum': 164, 'carry': 91}
        #10;
        $display("Test %0d: Inputs: a = 8'b10111011; b = 8'b01001100; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 164, 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011100; b = 8'b00110100; c = 8'b11100000; // Expected: {'sum': 72, 'carry': 180}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011100; b = 8'b00110100; c = 8'b11100000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 72, 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10001010; b = 8'b10000110; c = 8'b01010011; // Expected: {'sum': 95, 'carry': 130}
        #10;
        $display("Test %0d: Inputs: a = 8'b10001010; b = 8'b10000110; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 95, 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110011; b = 8'b01011100; c = 8'b11110001; // Expected: {'sum': 158, 'carry': 113}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110011; b = 8'b01011100; c = 8'b11110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 158, 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100001; b = 8'b00100000; c = 8'b01010011; // Expected: {'sum': 82, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100001; b = 8'b00100000; c = 8'b01010011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 82, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b01110100; c = 8'b00110000; // Expected: {'sum': 40, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b01110100; c = 8'b00110000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 40, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010100; b = 8'b10011111; c = 8'b00011111; // Expected: {'sum': 20, 'carry': 159}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010100; b = 8'b10011111; c = 8'b00011111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00111011; b = 8'b10011000; c = 8'b11111101; // Expected: {'sum': 94, 'carry': 185}
        #10;
        $display("Test %0d: Inputs: a = 8'b00111011; b = 8'b10011000; c = 8'b11111101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 94, 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101101; b = 8'b10100011; c = 8'b11000000; // Expected: {'sum': 142, 'carry': 225}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101101; b = 8'b10100011; c = 8'b11000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 142, 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00110111; b = 8'b00111101; c = 8'b01000100; // Expected: {'sum': 78, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b00110111; b = 8'b00111101; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 78, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11110010; b = 8'b00110001; c = 8'b11100100; // Expected: {'sum': 39, 'carry': 240}
        #10;
        $display("Test %0d: Inputs: a = 8'b11110010; b = 8'b00110001; c = 8'b11100100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 39, 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100100; b = 8'b00110001; c = 8'b10100010; // Expected: {'sum': 247, 'carry': 32}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100100; b = 8'b00110001; c = 8'b10100010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 247, 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101110; b = 8'b01010001; c = 8'b11000100; // Expected: {'sum': 59, 'carry': 196}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101110; b = 8'b01010001; c = 8'b11000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 59, 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001000; b = 8'b10010001; c = 8'b01000000; // Expected: {'sum': 25, 'carry': 192}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001000; b = 8'b10010001; c = 8'b01000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 25, 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11001001; b = 8'b00101000; c = 8'b00011000; // Expected: {'sum': 249, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 8'b11001001; b = 8'b00101000; c = 8'b00011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 249, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000110; b = 8'b00100001; c = 8'b10010001; // Expected: {'sum': 182, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000110; b = 8'b00100001; c = 8'b10010001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 182, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11000011; b = 8'b10000100; c = 8'b11111111; // Expected: {'sum': 184, 'carry': 199}
        #10;
        $display("Test %0d: Inputs: a = 8'b11000011; b = 8'b10000100; c = 8'b11111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 184, 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01010001; b = 8'b10111111; c = 8'b00110100; // Expected: {'sum': 218, 'carry': 53}
        #10;
        $display("Test %0d: Inputs: a = 8'b01010001; b = 8'b10111111; c = 8'b00110100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 218, 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11100100; b = 8'b01011010; c = 8'b10000010; // Expected: {'sum': 60, 'carry': 194}
        #10;
        $display("Test %0d: Inputs: a = 8'b11100100; b = 8'b01011010; c = 8'b10000010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 60, 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101001; b = 8'b01000011; c = 8'b11111001; // Expected: {'sum': 147, 'carry': 105}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101001; b = 8'b01000011; c = 8'b11111001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 147, 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00010111; b = 8'b10011010; c = 8'b01000100; // Expected: {'sum': 201, 'carry': 22}
        #10;
        $display("Test %0d: Inputs: a = 8'b00010111; b = 8'b10011010; c = 8'b01000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 201, 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101001; b = 8'b01100010; c = 8'b01000011; // Expected: {'sum': 200, 'carry': 99}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101001; b = 8'b01100010; c = 8'b01000011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 200, 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10010010; b = 8'b00011010; c = 8'b11111000; // Expected: {'sum': 112, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10010010; b = 8'b00011010; c = 8'b11111000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00000010; b = 8'b00111111; c = 8'b11000111; // Expected: {'sum': 250, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 8'b00000010; b = 8'b00111111; c = 8'b11000111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 250, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01100000; b = 8'b11110101; c = 8'b01110110; // Expected: {'sum': 227, 'carry': 116}
        #10;
        $display("Test %0d: Inputs: a = 8'b01100000; b = 8'b11110101; c = 8'b01110110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 227, 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111001; b = 8'b00111011; c = 8'b10111111; // Expected: {'sum': 253, 'carry': 59}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111001; b = 8'b00111011; c = 8'b10111111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 253, 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11101110; b = 8'b01110110; c = 8'b10011010; // Expected: {'sum': 2, 'carry': 254}
        #10;
        $display("Test %0d: Inputs: a = 8'b11101110; b = 8'b01110110; c = 8'b10011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000011; b = 8'b11000010; c = 8'b00101001; // Expected: {'sum': 168, 'carry': 67}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000011; b = 8'b11000010; c = 8'b00101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 168, 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101101; b = 8'b01000000; c = 8'b00110001; // Expected: {'sum': 220, 'carry': 33}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101101; b = 8'b01000000; c = 8'b00110001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 220, 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01111011; b = 8'b01000001; c = 8'b00101110; // Expected: {'sum': 20, 'carry': 107}
        #10;
        $display("Test %0d: Inputs: a = 8'b01111011; b = 8'b01000001; c = 8'b00101110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 20, 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10101000; b = 8'b01011101; c = 8'b01011000; // Expected: {'sum': 173, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b10101000; b = 8'b01011101; c = 8'b01011000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 173, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011001; b = 8'b10011010; c = 8'b01011010; // Expected: {'sum': 89, 'carry': 154}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011001; b = 8'b10011010; c = 8'b01011010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 89, 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01101100; b = 8'b00011110; c = 8'b11101001; // Expected: {'sum': 155, 'carry': 108}
        #10;
        $display("Test %0d: Inputs: a = 8'b01101100; b = 8'b00011110; c = 8'b11101001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 155, 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00100100; b = 8'b01011000; c = 8'b11011001; // Expected: {'sum': 165, 'carry': 88}
        #10;
        $display("Test %0d: Inputs: a = 8'b00100100; b = 8'b01011000; c = 8'b11011001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 165, 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b11011101; b = 8'b10101011; c = 8'b01000101; // Expected: {'sum': 51, 'carry': 205}
        #10;
        $display("Test %0d: Inputs: a = 8'b11011101; b = 8'b10101011; c = 8'b01000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 51, 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00011110; b = 8'b01110011; c = 8'b10111010; // Expected: {'sum': 215, 'carry': 58}
        #10;
        $display("Test %0d: Inputs: a = 8'b00011110; b = 8'b01110011; c = 8'b10111010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 215, 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101101; b = 8'b01101011; c = 8'b11110101; // Expected: {'sum': 179, 'carry': 109}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101101; b = 8'b01101011; c = 8'b11110101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 179, 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10011101; b = 8'b11111111; c = 8'b10000000; // Expected: {'sum': 226, 'carry': 157}
        #10;
        $display("Test %0d: Inputs: a = 8'b10011101; b = 8'b11111111; c = 8'b10000000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 226, 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b10100110; b = 8'b11001000; c = 8'b11110111; // Expected: {'sum': 153, 'carry': 230}
        #10;
        $display("Test %0d: Inputs: a = 8'b10100110; b = 8'b11001000; c = 8'b11110111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 153, 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b00101100; b = 8'b01101010; c = 8'b10000100; // Expected: {'sum': 194, 'carry': 44}
        #10;
        $display("Test %0d: Inputs: a = 8'b00101100; b = 8'b01101010; c = 8'b10000100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 194, 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 8'b01000101; b = 8'b11110000; c = 8'b11000101; // Expected: {'sum': 112, 'carry': 197}
        #10;
        $display("Test %0d: Inputs: a = 8'b01000101; b = 8'b11110000; c = 8'b11000101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 112, 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule