
`timescale 1ns / 1ps

module tb_N8_arithmetic_shifter;

    // Parameters
    
    parameter N = 8;
    
     
    // Inputs
    
    reg signed [7:0] data_in;
    
    reg  [2:0] shift_amount;
    
    reg   direction;
    
    
    // Outputs
    
    wire signed [7:0] data_out;
    
    
    // Instantiate the Unit Under Test (UUT)
    arithmetic_shifter  #( N ) uut (
        
        .data_in(data_in),
        
        .shift_amount(shift_amount),
        
        .direction(direction),
        
        
        .data_out(data_out)
        
    );

    // Clock generation 
    

    
    
    initial begin
        // Initialize Inputs
        
        data_in = 0;
        
        shift_amount = 0;
        
        direction = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 data_in = 8'b11111011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 0,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 4,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 5,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 6,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 7,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 8,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 9,
                 
                 data_out
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 10,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 11,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 12,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 13,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 14,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 15,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 16,
                 
                 data_out
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 17,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 206}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 18,
                 
                 data_out
                 , 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 19,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 20,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 21,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 22,
                 
                 data_out
                 , 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 23,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 24,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 25,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 26,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 27,
                 
                 data_out
                 , 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 28,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 29,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 30,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 31,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 32,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 33,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 34,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 35,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 36,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 37,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 38,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 39,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 40,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 41,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 42,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 43,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 44,
                 
                 data_out
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 45,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 46,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 47,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 48,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 49,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 50,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 51,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 52,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 53,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 54,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 55,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 56,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 57,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 58,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 59,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 60,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 119}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 61,
                 
                 data_out
                 , 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 62,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 63,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 64,
                 
                 data_out
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 65,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 66,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 67,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 68,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 69,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 70,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 71,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 72,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 73,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 74,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 75,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 76,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 77,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 78,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 79,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 80,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 81,
                 
                 data_out
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 82,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 83,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 206}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 84,
                 
                 data_out
                 , 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 85,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 86,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 89}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 87,
                 
                 data_out
                 , 
                 
                 89
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 88,
                 
                 data_out
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 89,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 90,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 91,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 92,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 93,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 94,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 133}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 95,
                 
                 data_out
                 , 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 96,
                 
                 data_out
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 97,
                 
                 data_out
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 98,
                 
                 data_out
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 99,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 100,
                 
                 data_out
                 , 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 101,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 102,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 103,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 104,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 105,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 106,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 107,
                 
                 data_out
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 108,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 109,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 110,
                 
                 data_out
                 , 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 111,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 112,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 113,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 203}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 114,
                 
                 data_out
                 , 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 115,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 116,
                 
                 data_out
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 117,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 118,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 119,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 120,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 121,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 122,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 123,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 124,
                 
                 data_out
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 125,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 126,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 127,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 173}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 128,
                 
                 data_out
                 , 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 129,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 130,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 131,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 132,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 133,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 134,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 135,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 136,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 137,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 138,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 139,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 140,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 141,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 142,
                 
                 data_out
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 143,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 144,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 145,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 146,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 147,
                 
                 data_out
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 148,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 149,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 150,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 151,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 152,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 153,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 154,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 155,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 156,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 157,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 158,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 159,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 160,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 161,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 162,
                 
                 data_out
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 163,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 164,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 165,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 166,
                 
                 data_out
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 167,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 168,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 169,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 170,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 171,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 172,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 173,
                 
                 data_out
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 174,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 175,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 176,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 177,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 178,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 179,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 180,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 181,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 182,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 183,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 184,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 185,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 186,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 187,
                 
                 data_out
                 , 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 188,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 211}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 189,
                 
                 data_out
                 , 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 190,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 191,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 192,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 193,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 194,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 195,
                 
                 data_out
                 , 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 196,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 197,
                 
                 data_out
                 , 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 198,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 199,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 200,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 201,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 202,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 94}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 203,
                 
                 data_out
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 204,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 205,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 206,
                 
                 data_out
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 207,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 208,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 191}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 209,
                 
                 data_out
                 , 
                 
                 191
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 210,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 211,
                 
                 data_out
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 212,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 213,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 223}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 214,
                 
                 data_out
                 , 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 215,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 216,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 217,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 218,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 219,
                 
                 data_out
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 91}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 220,
                 
                 data_out
                 , 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 221,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 222,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 223,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 224,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 225,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 226,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 227,
                 
                 data_out
                 , 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 228,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 229,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 230,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 231,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 232,
                 
                 data_out
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 233,
                 
                 data_out
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 234,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 235,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 236,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 237,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 238,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 83}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 239,
                 
                 data_out
                 , 
                 
                 83
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 240,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 241,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 242,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 243,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 244,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 245,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 246,
                 
                 data_out
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 247,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 248,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 249,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 250,
                 
                 data_out
                 , 
                 
                 131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 251,
                 
                 data_out
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 252,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 253,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 254,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 255,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 256,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 257,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 258,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 259,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 260,
                 
                 data_out
                 , 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 261,
                 
                 data_out
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 262,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 263,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 264,
                 
                 data_out
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 265,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 266,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 267,
                 
                 data_out
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 268,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 269,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 270,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 271,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 272,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 273,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 274,
                 
                 data_out
                 , 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 275,
                 
                 data_out
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 276,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 277,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 278,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 279,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 280,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 281,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 282,
                 
                 data_out
                 , 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 283,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 284,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 285,
                 
                 data_out
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 286,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 287,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 288,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 289,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 290,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 291,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 292,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 293,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 294,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 295,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 296,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 297,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 298,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 299,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 300,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 301,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 302,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 303,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 304,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 121}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 305,
                 
                 data_out
                 , 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 306,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 307,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 308,
                 
                 data_out
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 309,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 310,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 311,
                 
                 data_out
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 312,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 313,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 314,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 315,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 316,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 317,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 318,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 319,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 320,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 321,
                 
                 data_out
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 322,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 323,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 324,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 325,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 326,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 327,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 328,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 329,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 330,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 331,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 69}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 332,
                 
                 data_out
                 , 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 333,
                 
                 data_out
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 211}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 334,
                 
                 data_out
                 , 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 335,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 129}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 336,
                 
                 data_out
                 , 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 337,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 133}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 338,
                 
                 data_out
                 , 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 339,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 340,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 341,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 342,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 343,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 344,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 345,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 346,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 347,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 348,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 349,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 350,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 351,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 87}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 352,
                 
                 data_out
                 , 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 353,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 354,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 355,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 356,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 357,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 358,
                 
                 data_out
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 359,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 360,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 361,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 362,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 363,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 364,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 365,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 366,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 367,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 368,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 369,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 370,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 371,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 372,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 373,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 374,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 375,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 376,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 377,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 378,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 379,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 380,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 381,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 382,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 383,
                 
                 data_out
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 384,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 385,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 386,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 387,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 388,
                 
                 data_out
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 389,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 390,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 391,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 392,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 393,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 394,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 395,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 396,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 397,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 398,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 399,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 400,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 401,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 402,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 403,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 404,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 405,
                 
                 data_out
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 94}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 406,
                 
                 data_out
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 407,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 408,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 409,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 410,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 101}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 411,
                 
                 data_out
                 , 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 412,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 413,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 95}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 414,
                 
                 data_out
                 , 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 415,
                 
                 data_out
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 416,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 417,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 418,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 419,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 420,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 421,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 422,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 423,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 424,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 425,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 426,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 427,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 428,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 429,
                 
                 data_out
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 430,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 431,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 432,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 433,
                 
                 data_out
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 434,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 435,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 436,
                 
                 data_out
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 437,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 438,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 439,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 440,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 441,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 442,
                 
                 data_out
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 443,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 444,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 445,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 446,
                 
                 data_out
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 447,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 448,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 449,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 450,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 451,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 452,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 453,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 454,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 455,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 456,
                 
                 data_out
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 457,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 458,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 459,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 460,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 461,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 462,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 463,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 464,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 465,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 466,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 467,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 468,
                 
                 data_out
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 469,
                 
                 data_out
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 470,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 158}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 471,
                 
                 data_out
                 , 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 472,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 473,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 474,
                 
                 data_out
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 475,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 476,
                 
                 data_out
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 477,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 478,
                 
                 data_out
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 479,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 480,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 481,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 482,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 483,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 484,
                 
                 data_out
                 , 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 485,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 486,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 487,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 488,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 489,
                 
                 data_out
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 490,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 491,
                 
                 data_out
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 492,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 493,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 494,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 495,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 496,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 497,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 498,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 499,
                 
                 data_out
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 500,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 501,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 502,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 503,
                 
                 data_out
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 504,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 505,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 506,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 507,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 508,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 509,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 510,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 511,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 512,
                 
                 data_out
                 , 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 513,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 514,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 515,
                 
                 data_out
                 , 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 516,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 517,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 518,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 519,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 520,
                 
                 data_out
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 103}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 521,
                 
                 data_out
                 , 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 522,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 523,
                 
                 data_out
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 524,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 525,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 526,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 527,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 528,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 529,
                 
                 data_out
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 530,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 531,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 532,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 533,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 534,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 535,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 536,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 537,
                 
                 data_out
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 538,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 539,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 540,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 541,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 542,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 543,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 544,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 545,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 546,
                 
                 data_out
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 547,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 548,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 549,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 550,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 551,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 552,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 553,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 554,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 555,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 556,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 557,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 558,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 203}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 559,
                 
                 data_out
                 , 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 560,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 561,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 562,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 563,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 564,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 565,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 566,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 567,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 568,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 569,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 570,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 571,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 572,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 573,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 574,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 575,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 576,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 577,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 578,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 579,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 580,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 581,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 582,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 583,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 584,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 585,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 586,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 587,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 588,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 589,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 590,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 591,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 592,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 593,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 594,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 595,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 596,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 597,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 598,
                 
                 data_out
                 , 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 599,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 600,
                 
                 data_out
                 , 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 601,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 602,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 603,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 94}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 604,
                 
                 data_out
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 605,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 606,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 607,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 608,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 609,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 610,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 611,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 612,
                 
                 data_out
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 613,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 614,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 615,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 616,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 617,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 618,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 619,
                 
                 data_out
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 620,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 621,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 97}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 622,
                 
                 data_out
                 , 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 623,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 624,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 625,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 626,
                 
                 data_out
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 627,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 628,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 629,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 630,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 631,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 632,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 633,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 634,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 635,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 85}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 636,
                 
                 data_out
                 , 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 637,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 638,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 639,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 640,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 641,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 642,
                 
                 data_out
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 643,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 644,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 645,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 167}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 646,
                 
                 data_out
                 , 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 647,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 648,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 649,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 650,
                 
                 data_out
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 651,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 652,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 653,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 654,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 655,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 656,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 657,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 658,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 659,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 660,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 661,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 662,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 663,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 664,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 665,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 666,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 667,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 668,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 669,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 670,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 671,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 672,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 673,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 674,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 675,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 676,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 677,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 678,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 679,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 680,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 681,
                 
                 data_out
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 682,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 683,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 684,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 685,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 686,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 687,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 688,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 689,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 690,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 691,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 692,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 693,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 694,
                 
                 data_out
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 695,
                 
                 data_out
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 696,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 697,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 698,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 699,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 700,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 701,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 702,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 703,
                 
                 data_out
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 704,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 705,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 706,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 707,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 708,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 709,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 710,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 711,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 712,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 713,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 714,
                 
                 data_out
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 715,
                 
                 data_out
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 716,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 717,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 718,
                 
                 data_out
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 719,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 720,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 721,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 722,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 723,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 724,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 725,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 726,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 727,
                 
                 data_out
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 728,
                 
                 data_out
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 729,
                 
                 data_out
                 , 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 74}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 730,
                 
                 data_out
                 , 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 731,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 207}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 732,
                 
                 data_out
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 733,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 734,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 735,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 736,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 737,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 738,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 739,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 740,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 741,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 77}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 742,
                 
                 data_out
                 , 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 743,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 744,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 745,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 746,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 747,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 748,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 749,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 750,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 751,
                 
                 data_out
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 752,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 753,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 754,
                 
                 data_out
                 , 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 755,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 756,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 757,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 758,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 759,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 760,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 761,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 762,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 763,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 764,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 765,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 766,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 767,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 768,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 769,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 770,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 771,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 772,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 773,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 774,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 775,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 776,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 777,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 778,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 779,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 780,
                 
                 data_out
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 781,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 782,
                 
                 data_out
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 783,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 784,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 785,
                 
                 data_out
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 786,
                 
                 data_out
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 787,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 788,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 789,
                 
                 data_out
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 790,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 791,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 792,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 177}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 793,
                 
                 data_out
                 , 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 794,
                 
                 data_out
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 795,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 796,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 797,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 798,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 799,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 800,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 801,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 802,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 803,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 804,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 805,
                 
                 data_out
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 806,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 807,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 808,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 809,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 810,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 811,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 812,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 813,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 814,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 815,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 816,
                 
                 data_out
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 817,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 818,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 819,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 820,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 821,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 822,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 823,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 824,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 825,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 826,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 827,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 828,
                 
                 data_out
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 829,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 830,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 831,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 832,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 833,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 834,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 835,
                 
                 data_out
                 , 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 836,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 837,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 838,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 839,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 840,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 841,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 842,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 843,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 844,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 845,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 846,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 847,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 848,
                 
                 data_out
                 , 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 849,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 850,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 851,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 852,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 853,
                 
                 data_out
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 854,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 855,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 856,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 857,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 858,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 859,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 860,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 861,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 862,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 863,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 864,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 865,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 866,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 867,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 868,
                 
                 data_out
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 869,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 870,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 871,
                 
                 data_out
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 872,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 873,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 874,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 875,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 876,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 877,
                 
                 data_out
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 878,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 879,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 880,
                 
                 data_out
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 881,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 882,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 883,
                 
                 data_out
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 884,
                 
                 data_out
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 885,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 886,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 887,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 888,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 889,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 890,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 891,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 892,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 893,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 894,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 895,
                 
                 data_out
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 896,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 897,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 898,
                 
                 data_out
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 899,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 900,
                 
                 data_out
                 , 
                 
                 197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 901,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 902,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 903,
                 
                 data_out
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 904,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 905,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 906,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 907,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 137}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 908,
                 
                 data_out
                 , 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 909,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 910,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 911,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 912,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 913,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 914,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 915,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 916,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 917,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 918,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 919,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 920,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 921,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 922,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 923,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 924,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 925,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 926,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 927,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 928,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 929,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 930,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 931,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 932,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 933,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 934,
                 
                 data_out
                 , 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 935,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 936,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 937,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 938,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 939,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 940,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 941,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 942,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 943,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 944,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 945,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 946,
                 
                 data_out
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 947,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 103}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 948,
                 
                 data_out
                 , 
                 
                 103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 949,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 950,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 951,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 952,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 953,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 954,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 955,
                 
                 data_out
                 , 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 956,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 957,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 958,
                 
                 data_out
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 959,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 960,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 86}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 961,
                 
                 data_out
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 962,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 963,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 964,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 965,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 966,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 967,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 968,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 969,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 970,
                 
                 data_out
                 , 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 971,
                 
                 data_out
                 , 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 972,
                 
                 data_out
                 , 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 973,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 974,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 975,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 976,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 977,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 978,
                 
                 data_out
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 979,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 980,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 981,
                 
                 data_out
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 982,
                 
                 data_out
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 983,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 984,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 985,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 986,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 987,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 988,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 989,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 990,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 991,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 992,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 993,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 994,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 995,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 996,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 997,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 998,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 999,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1000,
                 
                 data_out
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1001,
                 
                 data_out
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1002,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1003,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1004,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1005,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1006,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1007,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1008,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1009,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1010,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1011,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1012,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1013,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1014,
                 
                 data_out
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1015,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1016,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1017,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1018,
                 
                 data_out
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1019,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1020,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1021,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1022,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1023,
                 
                 data_out
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1024,
                 
                 data_out
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1025,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1026,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1027,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1028,
                 
                 data_out
                 , 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1029,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1030,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 73}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1031,
                 
                 data_out
                 , 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 109}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1032,
                 
                 data_out
                 , 
                 
                 109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1033,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1034,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1035,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1036,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1037,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1038,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1039,
                 
                 data_out
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1040,
                 
                 data_out
                 , 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1041,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1042,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1043,
                 
                 data_out
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1044,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1045,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1046,
                 
                 data_out
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1047,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1048,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1049,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1050,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1051,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1052,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1053,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1054,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1055,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1056,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1057,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1058,
                 
                 data_out
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1059,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1060,
                 
                 data_out
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1061,
                 
                 data_out
                 , 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1062,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1063,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1064,
                 
                 data_out
                 , 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1065,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1066,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1067,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1068,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1069,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1070,
                 
                 data_out
                 , 
                 
                 115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1071,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1072,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1073,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1074,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1075,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1076,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1077,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1078,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1079,
                 
                 data_out
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1080,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1081,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1082,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1083,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1084,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1085,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1086,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1087,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1088,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1089,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1090,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1091,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1092,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1093,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1094,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1095,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1096,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1097,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1098,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1099,
                 
                 data_out
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1100,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1101,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1102,
                 
                 data_out
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1103,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1104,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1105,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1106,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1107,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1108,
                 
                 data_out
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1109,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1110,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1111,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1112,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1113,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1114,
                 
                 data_out
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1115,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1116,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1117,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1118,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1119,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1120,
                 
                 data_out
                 , 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1121,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1122,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1123,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1124,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1125,
                 
                 data_out
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1126,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1127,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1128,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1129,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1130,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1131,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1132,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1133,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1134,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 95}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1135,
                 
                 data_out
                 , 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1136,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1137,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1138,
                 
                 data_out
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1139,
                 
                 data_out
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1140,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1141,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1142,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1143,
                 
                 data_out
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1144,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1145,
                 
                 data_out
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1146,
                 
                 data_out
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1147,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1148,
                 
                 data_out
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1149,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1150,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1151,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1152,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1153,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1154,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1155,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1156,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1157,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1158,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1159,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1160,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1161,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1162,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1163,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1164,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1165,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1166,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1167,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1168,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1169,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1170,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1171,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1172,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1173,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1174,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1175,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1176,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1177,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1178,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1179,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1180,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1181,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1182,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1183,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1184,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1185,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 93}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1186,
                 
                 data_out
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1187,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1188,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1189,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1190,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1191,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 137}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1192,
                 
                 data_out
                 , 
                 
                 137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1193,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1194,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1195,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1196,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1197,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1198,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1199,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 158}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1200,
                 
                 data_out
                 , 
                 
                 158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1201,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1202,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1203,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1204,
                 
                 data_out
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1205,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1206,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1207,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1208,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1209,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1210,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1211,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1212,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1213,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1214,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1215,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1216,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1217,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1218,
                 
                 data_out
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1219,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1220,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1221,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1222,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1223,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1224,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1225,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1226,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1227,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1228,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1229,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1230,
                 
                 data_out
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1231,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1232,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1233,
                 
                 data_out
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 223}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1234,
                 
                 data_out
                 , 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1235,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1236,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1237,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1238,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1239,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1240,
                 
                 data_out
                 , 
                 
                 201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1241,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1242,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1243,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 177}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1244,
                 
                 data_out
                 , 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1245,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1246,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1247,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1248,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1249,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1250,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1251,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1252,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1253,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1254,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1255,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1256,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1257,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1258,
                 
                 data_out
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1259,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1260,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1261,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1262,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1263,
                 
                 data_out
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1264,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1265,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1266,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1267,
                 
                 data_out
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1268,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1269,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1270,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1271,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1272,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1273,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1274,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1275,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1276,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1277,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1278,
                 
                 data_out
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1279,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1280,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1281,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1282,
                 
                 data_out
                 , 
                 
                 233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1283,
                 
                 data_out
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1284,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1285,
                 
                 data_out
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1286,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1287,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1288,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1289,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1290,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1291,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1292,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1293,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1294,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1295,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1296,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1297,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1298,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1299,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1300,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1301,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1302,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1303,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1304,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1305,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1306,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1307,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 101}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1308,
                 
                 data_out
                 , 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1309,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1310,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1311,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1312,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1313,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1314,
                 
                 data_out
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1315,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1316,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 79}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1317,
                 
                 data_out
                 , 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1318,
                 
                 data_out
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1319,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1320,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1321,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1322,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1323,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1324,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1325,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1326,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1327,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1328,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1329,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1330,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1331,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1332,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1333,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1334,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1335,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1336,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1337,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1338,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1339,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1340,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1341,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1342,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1343,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1344,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1345,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1346,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1347,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1348,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1349,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1350,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1351,
                 
                 data_out
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1352,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1353,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1354,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1355,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1356,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1357,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1358,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1359,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1360,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1361,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1362,
                 
                 data_out
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1363,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1364,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1365,
                 
                 data_out
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1366,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1367,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1368,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1369,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1370,
                 
                 data_out
                 , 
                 
                 221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1371,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1372,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1373,
                 
                 data_out
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1374,
                 
                 data_out
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1375,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1376,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1377,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1378,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1379,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1380,
                 
                 data_out
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1381,
                 
                 data_out
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1382,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1383,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1384,
                 
                 data_out
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1385,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1386,
                 
                 data_out
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1387,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1388,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1389,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1390,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1391,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1392,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1393,
                 
                 data_out
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1394,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1395,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1396,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1397,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1398,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1399,
                 
                 data_out
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1400,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1401,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1402,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1403,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1404,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1405,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1406,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1407,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1408,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1409,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1410,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1411,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1412,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1413,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1414,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1415,
                 
                 data_out
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1416,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1417,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1418,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1419,
                 
                 data_out
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1420,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1421,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1422,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1423,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1424,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1425,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1426,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1427,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1428,
                 
                 data_out
                 , 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1429,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1430,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1431,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1432,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 147}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1433,
                 
                 data_out
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1434,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1435,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1436,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1437,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1438,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1439,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1440,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1441,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1442,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1443,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1444,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1445,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1446,
                 
                 data_out
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1447,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1448,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1449,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1450,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1451,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1452,
                 
                 data_out
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1453,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1454,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1455,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1456,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1457,
                 
                 data_out
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1458,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1459,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1460,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1461,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1462,
                 
                 data_out
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1463,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1464,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1465,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1466,
                 
                 data_out
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1467,
                 
                 data_out
                 , 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1468,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1469,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1470,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1471,
                 
                 data_out
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1472,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1473,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1474,
                 
                 data_out
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1475,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1476,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1477,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1478,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1479,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1480,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1481,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1482,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1483,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1484,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1485,
                 
                 data_out
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1486,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1487,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1488,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1489,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1490,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1491,
                 
                 data_out
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1492,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1493,
                 
                 data_out
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 117}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1494,
                 
                 data_out
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1495,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1496,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1497,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1498,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1499,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1500,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1501,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1502,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1503,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1504,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1505,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1506,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1507,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1508,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 229}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1509,
                 
                 data_out
                 , 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1510,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1511,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 65}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1512,
                 
                 data_out
                 , 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1513,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1514,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1515,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1516,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1517,
                 
                 data_out
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1518,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1519,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1520,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1521,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1522,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1523,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1524,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1525,
                 
                 data_out
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1526,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1527,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1528,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1529,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1530,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1531,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1532,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1533,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1534,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1535,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1536,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1537,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1538,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1539,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1540,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1541,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1542,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1543,
                 
                 data_out
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1544,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1545,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1546,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1547,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1548,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1549,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1550,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1551,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1552,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1553,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1554,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1555,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1556,
                 
                 data_out
                 , 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1557,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1558,
                 
                 data_out
                 , 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1559,
                 
                 data_out
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1560,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1561,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1562,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1563,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1564,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1565,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1566,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1567,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1568,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1569,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 194}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1570,
                 
                 data_out
                 , 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 141}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1571,
                 
                 data_out
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1572,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1573,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1574,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1575,
                 
                 data_out
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1576,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1577,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 181}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1578,
                 
                 data_out
                 , 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1579,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1580,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1581,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1582,
                 
                 data_out
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1583,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1584,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1585,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1586,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1587,
                 
                 data_out
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1588,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1589,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1590,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1591,
                 
                 data_out
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1592,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1593,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1594,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1595,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1596,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1597,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1598,
                 
                 data_out
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1599,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1600,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1601,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1602,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1603,
                 
                 data_out
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1604,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1605,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1606,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1607,
                 
                 data_out
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1608,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1609,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1610,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1611,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1612,
                 
                 data_out
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1613,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1614,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1615,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1616,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1617,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1618,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1619,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1620,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 79}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1621,
                 
                 data_out
                 , 
                 
                 79
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1622,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1623,
                 
                 data_out
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1624,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1625,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 203}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1626,
                 
                 data_out
                 , 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1627,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1628,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1629,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1630,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1631,
                 
                 data_out
                 , 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1632,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 194}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1633,
                 
                 data_out
                 , 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1634,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1635,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1636,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1637,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1638,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1639,
                 
                 data_out
                 , 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1640,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1641,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1642,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1643,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1644,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1645,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1646,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1647,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1648,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1649,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1650,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1651,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1652,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1653,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1654,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1655,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1656,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1657,
                 
                 data_out
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1658,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1659,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1660,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1661,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1662,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1663,
                 
                 data_out
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1664,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1665,
                 
                 data_out
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1666,
                 
                 data_out
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1667,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1668,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1669,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 143}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1670,
                 
                 data_out
                 , 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1671,
                 
                 data_out
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1672,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1673,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1674,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1675,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1676,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1677,
                 
                 data_out
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1678,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1679,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1680,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1681,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1682,
                 
                 data_out
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1683,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1684,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1685,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1686,
                 
                 data_out
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1687,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1688,
                 
                 data_out
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1689,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1690,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1691,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1692,
                 
                 data_out
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1693,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1694,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1695,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1696,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 229}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1697,
                 
                 data_out
                 , 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1698,
                 
                 data_out
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1699,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1700,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1701,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1702,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1703,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1704,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1705,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1706,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1707,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1708,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1709,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1710,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1711,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1712,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1713,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1714,
                 
                 data_out
                 , 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1715,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1716,
                 
                 data_out
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1717,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1718,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1719,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1720,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1721,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1722,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1723,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1724,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1725,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1726,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1727,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1728,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1729,
                 
                 data_out
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1730,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1731,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1732,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1733,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1734,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1735,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1736,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1737,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1738,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1739,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1740,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1741,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 127}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1742,
                 
                 data_out
                 , 
                 
                 127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1743,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1744,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1745,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1746,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1747,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1748,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1749,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1750,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1751,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1752,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1753,
                 
                 data_out
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1754,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1755,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1756,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1757,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1758,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1759,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1760,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1761,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1762,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1763,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1764,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1765,
                 
                 data_out
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1766,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1767,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1768,
                 
                 data_out
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1769,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1770,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1771,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1772,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1773,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1774,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1775,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1776,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1777,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1778,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1779,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1780,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1781,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1782,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1783,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1784,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1785,
                 
                 data_out
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1786,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1787,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1788,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1789,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1790,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1791,
                 
                 data_out
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1792,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1793,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1794,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1795,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1796,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1797,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1798,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1799,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1800,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1801,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1802,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1803,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1804,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1805,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1806,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1807,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1808,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1809,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1810,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1811,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1812,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1813,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1814,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1815,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1816,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1817,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 211}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1818,
                 
                 data_out
                 , 
                 
                 211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1819,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1820,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1821,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1822,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1823,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1824,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1825,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 123}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1826,
                 
                 data_out
                 , 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1827,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1828,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 223}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1829,
                 
                 data_out
                 , 
                 
                 223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1830,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1831,
                 
                 data_out
                 , 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1832,
                 
                 data_out
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1833,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1834,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1835,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1836,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1837,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1838,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1839,
                 
                 data_out
                 , 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1840,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1841,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1842,
                 
                 data_out
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1843,
                 
                 data_out
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1844,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1845,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1846,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1847,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1848,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1849,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1850,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1851,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1852,
                 
                 data_out
                 , 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1853,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1854,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1855,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1856,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1857,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1858,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1859,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1860,
                 
                 data_out
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1861,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1862,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1863,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1864,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1865,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1866,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1867,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1868,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1869,
                 
                 data_out
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1870,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1871,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1872,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1873,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1874,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1875,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1876,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1877,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1878,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1879,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1880,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1881,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1882,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1883,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1884,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1885,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1886,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1887,
                 
                 data_out
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1888,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1889,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1890,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1891,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1892,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1893,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1894,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1895,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1896,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1897,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1898,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1899,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1900,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1901,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1902,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1903,
                 
                 data_out
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1904,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1905,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1906,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1907,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1908,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1909,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1910,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1911,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1912,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1913,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1914,
                 
                 data_out
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1915,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1916,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1917,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1918,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1919,
                 
                 data_out
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1920,
                 
                 data_out
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1921,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1922,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1923,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1924,
                 
                 data_out
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1925,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1926,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1927,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1928,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 139}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1929,
                 
                 data_out
                 , 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 151}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1930,
                 
                 data_out
                 , 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1931,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1932,
                 
                 data_out
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1933,
                 
                 data_out
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1934,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1935,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1936,
                 
                 data_out
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1937,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1938,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1939,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1940,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1941,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1942,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1943,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1944,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1945,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1946,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1947,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1948,
                 
                 data_out
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1949,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1950,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1951,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1952,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 194}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1953,
                 
                 data_out
                 , 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1954,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1955,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1956,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1957,
                 
                 data_out
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1958,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1959,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1960,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1961,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1962,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1963,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1964,
                 
                 data_out
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1965,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1966,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1967,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1968,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1969,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1970,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1971,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1972,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1973,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1974,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1975,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1976,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1977,
                 
                 data_out
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1978,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1979,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1980,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1981,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1982,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1983,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1984,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1985,
                 
                 data_out
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1986,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1987,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1988,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1989,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1990,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1991,
                 
                 data_out
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1992,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1993,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1994,
                 
                 data_out
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1995,
                 
                 data_out
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1996,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 1997,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1998,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 1999,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2000,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2001,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2002,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2003,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2004,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2005,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2006,
                 
                 data_out
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2007,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2008,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2009,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2010,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2011,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2012,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2013,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2014,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2015,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2016,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2017,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2018,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2019,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2020,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2021,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2022,
                 
                 data_out
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2023,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2024,
                 
                 data_out
                 , 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2025,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2026,
                 
                 data_out
                 , 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2027,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2028,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2029,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2030,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2031,
                 
                 data_out
                 , 
                 
                 235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2032,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2033,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2034,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2035,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2036,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2037,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2038,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2039,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2040,
                 
                 data_out
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2041,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2042,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2043,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 111}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2044,
                 
                 data_out
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2045,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2046,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2047,
                 
                 data_out
                 , 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2048,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2049,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2050,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2051,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2052,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2053,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2054,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2055,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2056,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2057,
                 
                 data_out
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2058,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2059,
                 
                 data_out
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2060,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2061,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2062,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2063,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2064,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2065,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2066,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2067,
                 
                 data_out
                 , 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2068,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2069,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2070,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2071,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2072,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2073,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2074,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2075,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2076,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2077,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2078,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2079,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2080,
                 
                 data_out
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2081,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2082,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2083,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2084,
                 
                 data_out
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2085,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2086,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 194}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2087,
                 
                 data_out
                 , 
                 
                 194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2088,
                 
                 data_out
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2089,
                 
                 data_out
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2090,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2091,
                 
                 data_out
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2092,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2093,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2094,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2095,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2096,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2097,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2098,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2099,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2100,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2101,
                 
                 data_out
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2102,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2103,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2104,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2105,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2106,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2107,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2108,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2109,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2110,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2111,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2112,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2113,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2114,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2115,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2116,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2117,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2118,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2119,
                 
                 data_out
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2120,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2121,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2122,
                 
                 data_out
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2123,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2124,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2125,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2126,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2127,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2128,
                 
                 data_out
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2129,
                 
                 data_out
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2130,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2131,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 73}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2132,
                 
                 data_out
                 , 
                 
                 73
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2133,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2134,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2135,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2136,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2137,
                 
                 data_out
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2138,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2139,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2140,
                 
                 data_out
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2141,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2142,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2143,
                 
                 data_out
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2144,
                 
                 data_out
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2145,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2146,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2147,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 149}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2148,
                 
                 data_out
                 , 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2149,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2150,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2151,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2152,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2153,
                 
                 data_out
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2154,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2155,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2156,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2157,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2158,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2159,
                 
                 data_out
                 , 
                 
                 213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2160,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2161,
                 
                 data_out
                 , 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2162,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2163,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2164,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2165,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2166,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 167}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2167,
                 
                 data_out
                 , 
                 
                 167
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2168,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2169,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2170,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2171,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2172,
                 
                 data_out
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2173,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2174,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2175,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2176,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 123}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2177,
                 
                 data_out
                 , 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2178,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2179,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2180,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2181,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2182,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2183,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2184,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2185,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2186,
                 
                 data_out
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2187,
                 
                 data_out
                 , 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2188,
                 
                 data_out
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2189,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2190,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2191,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2192,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2193,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2194,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2195,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2196,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2197,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2198,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 93}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2199,
                 
                 data_out
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2200,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2201,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2202,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2203,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2204,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2205,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2206,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2207,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2208,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 74}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2209,
                 
                 data_out
                 , 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2210,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2211,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2212,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 157}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2213,
                 
                 data_out
                 , 
                 
                 157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2214,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2215,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 161}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2216,
                 
                 data_out
                 , 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2217,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2218,
                 
                 data_out
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2219,
                 
                 data_out
                 , 
                 
                 166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2220,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2221,
                 
                 data_out
                 , 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2222,
                 
                 data_out
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2223,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2224,
                 
                 data_out
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2225,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2226,
                 
                 data_out
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2227,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2228,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2229,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2230,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2231,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2232,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2233,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2234,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2235,
                 
                 data_out
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2236,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2237,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2238,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2239,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2240,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 111}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2241,
                 
                 data_out
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2242,
                 
                 data_out
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 91}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2243,
                 
                 data_out
                 , 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2244,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2245,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2246,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2247,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2248,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2249,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2250,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2251,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2252,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2253,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2254,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2255,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2256,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2257,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2258,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2259,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2260,
                 
                 data_out
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2261,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2262,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2263,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2264,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2265,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2266,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2267,
                 
                 data_out
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2268,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2269,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2270,
                 
                 data_out
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2271,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2272,
                 
                 data_out
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2273,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2274,
                 
                 data_out
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2275,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2276,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2277,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 173}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2278,
                 
                 data_out
                 , 
                 
                 173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2279,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2280,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2281,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2282,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2283,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 163}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2284,
                 
                 data_out
                 , 
                 
                 163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2285,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2286,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2287,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2288,
                 
                 data_out
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2289,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2290,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2291,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2292,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2293,
                 
                 data_out
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2294,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2295,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2296,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2297,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2298,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2299,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2300,
                 
                 data_out
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2301,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2302,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2303,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2304,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2305,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2306,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2307,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2308,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2309,
                 
                 data_out
                 , 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2310,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 229}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2311,
                 
                 data_out
                 , 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2312,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2313,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2314,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2315,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2316,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2317,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2318,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2319,
                 
                 data_out
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2320,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2321,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2322,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2323,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2324,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2325,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2326,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2327,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2328,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2329,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2330,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2331,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2332,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2333,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2334,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2335,
                 
                 data_out
                 , 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2336,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2337,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2338,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2339,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2340,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2341,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2342,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2343,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2344,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2345,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2346,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2347,
                 
                 data_out
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2348,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2349,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2350,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2351,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2352,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2353,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2354,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2355,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2356,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2357,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2358,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2359,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2360,
                 
                 data_out
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2361,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2362,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2363,
                 
                 data_out
                 , 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2364,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2365,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2366,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2367,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2368,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2369,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2370,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2371,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2372,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2373,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2374,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2375,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2376,
                 
                 data_out
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2377,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2378,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2379,
                 
                 data_out
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2380,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2381,
                 
                 data_out
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2382,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2383,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2384,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2385,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2386,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2387,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2388,
                 
                 data_out
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2389,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2390,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2391,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2392,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2393,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2394,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2395,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2396,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2397,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2398,
                 
                 data_out
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2399,
                 
                 data_out
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2400,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2401,
                 
                 data_out
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2402,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2403,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2404,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2405,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2406,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2407,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2408,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2409,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2410,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2411,
                 
                 data_out
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2412,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2413,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2414,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2415,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2416,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2417,
                 
                 data_out
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2418,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2419,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2420,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2421,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2422,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2423,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2424,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2425,
                 
                 data_out
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2426,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2427,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2428,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2429,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2430,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2431,
                 
                 data_out
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2432,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2433,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2434,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2435,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2436,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2437,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2438,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2439,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2440,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2441,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2442,
                 
                 data_out
                 , 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2443,
                 
                 data_out
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2444,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2445,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2446,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2447,
                 
                 data_out
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2448,
                 
                 data_out
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2449,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2450,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2451,
                 
                 data_out
                 , 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2452,
                 
                 data_out
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 181}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2453,
                 
                 data_out
                 , 
                 
                 181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2454,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2455,
                 
                 data_out
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2456,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2457,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2458,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2459,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2460,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2461,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2462,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2463,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2464,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2465,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2466,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2467,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2468,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2469,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2470,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2471,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2472,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2473,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2474,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2475,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2476,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2477,
                 
                 data_out
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2478,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2479,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2480,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2481,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2482,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2483,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2484,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2485,
                 
                 data_out
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2486,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2487,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2488,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2489,
                 
                 data_out
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2490,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2491,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2492,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2493,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2494,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2495,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2496,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2497,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2498,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2499,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2500,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2501,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2502,
                 
                 data_out
                 , 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2503,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2504,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2505,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2506,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2507,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2508,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2509,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2510,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2511,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2512,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2513,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2514,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2515,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2516,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2517,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2518,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2519,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2520,
                 
                 data_out
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2521,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2522,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2523,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2524,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2525,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2526,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2527,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2528,
                 
                 data_out
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2529,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2530,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2531,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2532,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101100; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101100; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2533,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2534,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2535,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2536,
                 
                 data_out
                 , 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2537,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2538,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2539,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2540,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2541,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 59}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2542,
                 
                 data_out
                 , 
                 
                 59
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2543,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2544,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2545,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2546,
                 
                 data_out
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2547,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2548,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2549,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2550,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2551,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2552,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2553,
                 
                 data_out
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2554,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2555,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2556,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2557,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2558,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2559,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 206}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2560,
                 
                 data_out
                 , 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2561,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2562,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 229}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2563,
                 
                 data_out
                 , 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2564,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2565,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2566,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2567,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2568,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2569,
                 
                 data_out
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2570,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2571,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2572,
                 
                 data_out
                 , 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2573,
                 
                 data_out
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2574,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2575,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2576,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2577,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2578,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2579,
                 
                 data_out
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2580,
                 
                 data_out
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2581,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2582,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2583,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2584,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2585,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2586,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2587,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2588,
                 
                 data_out
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2589,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2590,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 86}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2591,
                 
                 data_out
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2592,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2593,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2594,
                 
                 data_out
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2595,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2596,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2597,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2598,
                 
                 data_out
                 , 
                 
                 214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2599,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2600,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2601,
                 
                 data_out
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2602,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2603,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2604,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2605,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2606,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2607,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2608,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2609,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2610,
                 
                 data_out
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2611,
                 
                 data_out
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2612,
                 
                 data_out
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2613,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2614,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2615,
                 
                 data_out
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2616,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2617,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2618,
                 
                 data_out
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 21}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2619,
                 
                 data_out
                 , 
                 
                 21
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2620,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 151}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2621,
                 
                 data_out
                 , 
                 
                 151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2622,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2623,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2624,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2625,
                 
                 data_out
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2626,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2627,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2628,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 37}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2629,
                 
                 data_out
                 , 
                 
                 37
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2630,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2631,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2632,
                 
                 data_out
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2633,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2634,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2635,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2636,
                 
                 data_out
                 , 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2637,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2638,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2639,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2640,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2641,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2642,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2643,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2644,
                 
                 data_out
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2645,
                 
                 data_out
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2646,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2647,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2648,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2649,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2650,
                 
                 data_out
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2651,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2652,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2653,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2654,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2655,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2656,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2657,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2658,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2659,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2660,
                 
                 data_out
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2661,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 94}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2662,
                 
                 data_out
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2663,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2664,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2665,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2666,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2667,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2668,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2669,
                 
                 data_out
                 , 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2670,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2671,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2672,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2673,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2674,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2675,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2676,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2677,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 179}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2678,
                 
                 data_out
                 , 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2679,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2680,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2681,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2682,
                 
                 data_out
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2683,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2684,
                 
                 data_out
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2685,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2686,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2687,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2688,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2689,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2690,
                 
                 data_out
                 , 
                 
                 178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2691,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2692,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2693,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2694,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2695,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2696,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2697,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2698,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2699,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2700,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2701,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2702,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2703,
                 
                 data_out
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 67}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2704,
                 
                 data_out
                 , 
                 
                 67
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2705,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2706,
                 
                 data_out
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 202}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2707,
                 
                 data_out
                 , 
                 
                 202
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2708,
                 
                 data_out
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2709,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 179}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2710,
                 
                 data_out
                 , 
                 
                 179
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2711,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2712,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2713,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2714,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2715,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2716,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2717,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2718,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2719,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2720,
                 
                 data_out
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2721,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2722,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2723,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 141}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2724,
                 
                 data_out
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2725,
                 
                 data_out
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2726,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2727,
                 
                 data_out
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2728,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2729,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2730,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2731,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2732,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2733,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2734,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2735,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2736,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2737,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2738,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2739,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2740,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2741,
                 
                 data_out
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2742,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2743,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2744,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2745,
                 
                 data_out
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2746,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2747,
                 
                 data_out
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2748,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2749,
                 
                 data_out
                 , 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2750,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2751,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2752,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2753,
                 
                 data_out
                 , 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2754,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2755,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2756,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2757,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2758,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2759,
                 
                 data_out
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2760,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101100; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101100; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2761,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2762,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2763,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2764,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2765,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2766,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2767,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2768,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2769,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2770,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2771,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2772,
                 
                 data_out
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001110; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001110; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2773,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2774,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2775,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2776,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2777,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2778,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2779,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2780,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2781,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2782,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2783,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2784,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2785,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2786,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2787,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2788,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2789,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2790,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2791,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2792,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2793,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2794,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2795,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2796,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2797,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2798,
                 
                 data_out
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2799,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2800,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2801,
                 
                 data_out
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2802,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2803,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 149}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2804,
                 
                 data_out
                 , 
                 
                 149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2805,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2806,
                 
                 data_out
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2807,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2808,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2809,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2810,
                 
                 data_out
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2811,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2812,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2813,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2814,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2815,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2816,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2817,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2818,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2819,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2820,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2821,
                 
                 data_out
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2822,
                 
                 data_out
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2823,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2824,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2825,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2826,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2827,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2828,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2829,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2830,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2831,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2832,
                 
                 data_out
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2833,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2834,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2835,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2836,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101001; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101001; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2837,
                 
                 data_out
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2838,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2839,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2840,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2841,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2842,
                 
                 data_out
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2843,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2844,
                 
                 data_out
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2845,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2846,
                 
                 data_out
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2847,
                 
                 data_out
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2848,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2849,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2850,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2851,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2852,
                 
                 data_out
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2853,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2854,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2855,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2856,
                 
                 data_out
                 , 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2857,
                 
                 data_out
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2858,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2859,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2860,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2861,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2862,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2863,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2864,
                 
                 data_out
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2865,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2866,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2867,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2868,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2869,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2870,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 139}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2871,
                 
                 data_out
                 , 
                 
                 139
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2872,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000000; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000000; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2873,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2874,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 4}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2875,
                 
                 data_out
                 , 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2876,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2877,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2878,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2879,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2880,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2881,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2882,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011111; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011111; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2883,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2884,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2885,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2886,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2887,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2888,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2889,
                 
                 data_out
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2890,
                 
                 data_out
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2891,
                 
                 data_out
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2892,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2893,
                 
                 data_out
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2894,
                 
                 data_out
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2895,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2896,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2897,
                 
                 data_out
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2898,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2899,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2900,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2901,
                 
                 data_out
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2902,
                 
                 data_out
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2903,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2904,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2905,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2906,
                 
                 data_out
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100111; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100111; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2907,
                 
                 data_out
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2908,
                 
                 data_out
                 , 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2909,
                 
                 data_out
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2910,
                 
                 data_out
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2911,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2912,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2913,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2914,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2915,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2916,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2917,
                 
                 data_out
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2918,
                 
                 data_out
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2919,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2920,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2921,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2922,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2923,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2924,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2925,
                 
                 data_out
                 , 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010101; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010101; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2926,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2927,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 227}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2928,
                 
                 data_out
                 , 
                 
                 227
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001011; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001011; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2929,
                 
                 data_out
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2930,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2931,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2932,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2933,
                 
                 data_out
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2934,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2935,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2936,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2937,
                 
                 data_out
                 , 
                 
                 113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011111; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011111; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2938,
                 
                 data_out
                 , 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2939,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2940,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2941,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2942,
                 
                 data_out
                 , 
                 
                 199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2943,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2944,
                 
                 data_out
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2945,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2946,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2947,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2948,
                 
                 data_out
                 , 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2949,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110111; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110111; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2950,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2951,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2952,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2953,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111110; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111110; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2954,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011000; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011000; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2955,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2956,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2957,
                 
                 data_out
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2958,
                 
                 data_out
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2959,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110011; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110011; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2960,
                 
                 data_out
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2961,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100001; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100001; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2962,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2963,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2964,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2965,
                 
                 data_out
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2966,
                 
                 data_out
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2967,
                 
                 data_out
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2968,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2969,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11011000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11011000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2970,
                 
                 data_out
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2971,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2972,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2973,
                 
                 data_out
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2974,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2975,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2976,
                 
                 data_out
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2977,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2978,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2979,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2980,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2981,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2982,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2983,
                 
                 data_out
                 , 
                 
                 241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2984,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2985,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2986,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 206}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2987,
                 
                 data_out
                 , 
                 
                 206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2988,
                 
                 data_out
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2989,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2990,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001100; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001100; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2991,
                 
                 data_out
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000010; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000010; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2992,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100011; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100011; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2993,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2994,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2995,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2996,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001000; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001000; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2997,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 2998,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010111; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010111; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 2999,
                 
                 data_out
                 , 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3000,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3001,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3002,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 193}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3003,
                 
                 data_out
                 , 
                 
                 193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3004,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3005,
                 
                 data_out
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3006,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3007,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3008,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111010; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111010; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3009,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3010,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3011,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 77}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3012,
                 
                 data_out
                 , 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001111; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001111; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3013,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110101; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110101; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3014,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3015,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3016,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3017,
                 
                 data_out
                 , 
                 
                 239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010001; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010001; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3018,
                 
                 data_out
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001101; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001101; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3019,
                 
                 data_out
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010011; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010011; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3020,
                 
                 data_out
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3021,
                 
                 data_out
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3022,
                 
                 data_out
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3023,
                 
                 data_out
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3024,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111001; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111001; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3025,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00000111; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00000111; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3026,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11010001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11010001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3027,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010101; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010101; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3028,
                 
                 data_out
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101110; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101110; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3029,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011001; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 153}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011001; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3030,
                 
                 data_out
                 , 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3031,
                 
                 data_out
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3032,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3033,
                 
                 data_out
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110100; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110100; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3034,
                 
                 data_out
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100111; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100111; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3035,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3036,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101111; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101111; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3037,
                 
                 data_out
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100001; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100001; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3038,
                 
                 data_out
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3039,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101000; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101000; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3040,
                 
                 data_out
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111011; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111011; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3041,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3042,
                 
                 data_out
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3043,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3044,
                 
                 data_out
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3045,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111010; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111010; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3046,
                 
                 data_out
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111001; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111001; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3047,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00011101; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00011101; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3048,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11110010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11110010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3049,
                 
                 data_out
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111110; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111110; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3050,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3051,
                 
                 data_out
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3052,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3053,
                 
                 data_out
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3054,
                 
                 data_out
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001100; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001100; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3055,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3056,
                 
                 data_out
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3057,
                 
                 data_out
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110000; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110000; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3058,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001011; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001011; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3059,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110010; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110010; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3060,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11001111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11001111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3061,
                 
                 data_out
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3062,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3063,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3064,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110010; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110010; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3065,
                 
                 data_out
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100011; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 99}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100011; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3066,
                 
                 data_out
                 , 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3067,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011100; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011100; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3068,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110111; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110111; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3069,
                 
                 data_out
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110011; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110011; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3070,
                 
                 data_out
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3071,
                 
                 data_out
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3072,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111111; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111111; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3073,
                 
                 data_out
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01100010; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01100010; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3074,
                 
                 data_out
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010000; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010000; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3075,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00110101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00110101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3076,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3077,
                 
                 data_out
                 , 
                 
                 254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000001; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 65}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000001; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3078,
                 
                 data_out
                 , 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11111001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11111001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3079,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001110; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001110; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3080,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b100; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b100; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3081,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b000; direction = 1'b0; // Expected: {'data_out': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b000; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3082,
                 
                 data_out
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00001010; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00001010; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3083,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3084,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01011010; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01011010; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3085,
                 
                 data_out
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3086,
                 
                 data_out
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3087,
                 
                 data_out
                 , 
                 
                 226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101101; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101101; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3088,
                 
                 data_out
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111111; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111111; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3089,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101101; shift_amount = 3'b110; direction = 1'b0; // Expected: {'data_out': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101101; shift_amount = 3'b110; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3090,
                 
                 data_out
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01110111; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 1}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01110111; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3091,
                 
                 data_out
                 , 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010110; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010110; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3092,
                 
                 data_out
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10101010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10101010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3093,
                 
                 data_out
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01111101; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01111101; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3094,
                 
                 data_out
                 , 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10100000; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10100000; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3095,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01010011; shift_amount = 3'b101; direction = 1'b1; // Expected: {'data_out': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01010011; shift_amount = 3'b101; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3096,
                 
                 data_out
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10011101; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10011101; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3097,
                 
                 data_out
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010000; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010000; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3098,
                 
                 data_out
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001101; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001101; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3099,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110010; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110010; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3100,
                 
                 data_out
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10001110; shift_amount = 3'b000; direction = 1'b1; // Expected: {'data_out': 142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10001110; shift_amount = 3'b000; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3101,
                 
                 data_out
                 , 
                 
                 142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01001001; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01001001; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3102,
                 
                 data_out
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100110; shift_amount = 3'b110; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100110; shift_amount = 3'b110; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3103,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010111; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 229}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010111; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3104,
                 
                 data_out
                 , 
                 
                 229
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00100100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00100100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3105,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101110; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101110; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3106,
                 
                 data_out
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11100010; shift_amount = 3'b011; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11100010; shift_amount = 3'b011; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3107,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111101; shift_amount = 3'b101; direction = 1'b0; // Expected: {'data_out': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111101; shift_amount = 3'b101; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3108,
                 
                 data_out
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10010001; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10010001; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3109,
                 
                 data_out
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101100; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101100; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3110,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10110011; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10110011; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3111,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00010001; shift_amount = 3'b011; direction = 1'b0; // Expected: {'data_out': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00010001; shift_amount = 3'b011; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3112,
                 
                 data_out
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00111100; shift_amount = 3'b001; direction = 1'b1; // Expected: {'data_out': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00111100; shift_amount = 3'b001; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3113,
                 
                 data_out
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10000100; shift_amount = 3'b001; direction = 1'b0; // Expected: {'data_out': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10000100; shift_amount = 3'b001; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3114,
                 
                 data_out
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101111; shift_amount = 3'b111; direction = 1'b0; // Expected: {'data_out': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101111; shift_amount = 3'b111; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3115,
                 
                 data_out
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b10111110; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b10111110; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3116,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11101110; shift_amount = 3'b010; direction = 1'b1; // Expected: {'data_out': 251}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11101110; shift_amount = 3'b010; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3117,
                 
                 data_out
                 , 
                 
                 251
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01101101; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01101101; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3118,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b11000000; shift_amount = 3'b100; direction = 1'b1; // Expected: {'data_out': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b11000000; shift_amount = 3'b100; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3119,
                 
                 data_out
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b01000100; shift_amount = 3'b111; direction = 1'b1; // Expected: {'data_out': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b01000100; shift_amount = 3'b111; direction = 1'b1; | Outputs: data_out=%b | Expected: data_out=%d",
                 3120,
                 
                 data_out
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 data_in = 8'b00101011; shift_amount = 3'b010; direction = 1'b0; // Expected: {'data_out': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: data_in = 8'b00101011; shift_amount = 3'b010; direction = 1'b0; | Outputs: data_out=%b | Expected: data_out=%d",
                 3121,
                 
                 data_out
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule