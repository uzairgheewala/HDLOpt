
`timescale 1ns / 1ps

module tb_N4_carry_save_adder_l2;

    // Parameters
    
    parameter N = 4;
    
     
    // Inputs
    
    reg  [3:0] a;
    
    reg  [3:0] b;
    
    reg  [3:0] c;
    
    
    // Outputs
    
    wire  [3:0] sum;
    
    wire  [3:0] carry;
    
    
    // Instantiate the Unit Under Test (UUT)
    carry_save_adder_l2  #( N ) uut (
        
        .a(a),
        
        .b(b),
        
        .c(c),
        
        
        .sum(sum),
        
        .carry(carry)
        
    );
    
    initial begin
        // Initialize Inputs
        
        a = 0;
        
        b = 0;
        
        c = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        a = 4'b1000; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 0,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 4,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 5,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 6,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 7,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 8,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 9,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 10,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 11,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 12,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 13,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 14,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 5, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 15,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 16,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 17,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 18,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 19,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 20,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 21,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 22,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 23,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 24,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 25,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 26,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 27,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 28,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 29,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 30,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 31,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 32,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 33,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 34,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 35,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 36,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 37,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 38,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 39,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 40,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 41,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 42,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 43,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 44,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 45,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 46,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 47,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 7, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 48,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 49,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 50,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 51,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 52,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 53,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 54,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 55,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 56,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 57,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 58,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 59,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 60,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 5, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 61,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 62,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 63,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 64,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 65,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 66,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 67,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 68,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 69,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 70,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 71,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 72,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 73,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 74,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 75,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 76,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 77,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 78,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 79,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 80,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 81,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 82,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 83,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 84,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 85,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 86,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 87,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 88,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 89,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 90,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 91,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 92,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 93,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 94,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 13, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 95,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 96,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 97,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 98,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 99,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 6, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 12, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 0, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 2, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 8, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 1, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 4, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 13, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 1, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 7, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 5, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 13, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 6, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 3, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 0, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 14, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 10, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 5, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 6, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 9, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 3, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 8, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 3, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 9, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 12, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 12, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 9, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 4, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 10, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 14, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 10, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 1, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 10, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 14, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 5, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 2, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 9, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 3, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 663,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 0, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 664,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 665,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 666,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 3, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 667,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 668,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 669,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 670,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 671,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 672,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 673,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 674,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 675,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 676,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 677,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 678,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 679,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 680,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 681,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 682,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 683,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 684,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 685,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 686,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 687,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 688,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 689,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 690,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 691,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 14, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 692,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 693,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 694,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 695,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 696,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 697,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 698,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 699,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 700,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 701,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 702,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 703,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 704,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 705,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 706,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 707,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 708,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 709,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 710,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 711,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 712,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 713,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 714,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 715,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 716,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 8, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 717,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 718,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 719,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 720,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 721,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 722,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 723,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 724,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 725,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 726,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 727,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 728,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 729,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 730,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 731,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 732,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 733,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 734,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 735,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 736,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 737,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 738,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 739,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 740,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 741,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 742,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 743,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 744,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 745,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 746,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 747,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 748,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 2, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 749,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 750,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 751,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 752,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 753,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 754,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 755,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 756,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 757,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 758,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 759,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 760,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 761,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 762,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 763,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 764,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 765,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 766,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 767,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 768,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 769,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 770,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 0, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 771,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 772,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 773,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 774,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 775,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 776,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 777,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 778,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 11, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 779,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 780,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 781,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 782,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 783,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 784,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 785,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 0, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 786,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 787,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 788,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 789,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 790,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 791,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 792,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 793,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 794,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 795,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 796,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 797,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 798,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 799,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 800,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 801,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 802,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 803,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 804,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 9, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 805,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 806,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 807,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 808,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 10, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 809,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 810,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 811,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 812,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 813,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 814,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 14, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 815,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 816,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 817,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 818,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 819,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 820,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 821,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 822,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 823,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 824,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 825,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 826,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 827,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 828,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 829,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 830,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 831,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 832,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 833,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 834,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 835,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 836,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 837,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 838,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 839,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 840,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 841,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 842,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 843,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 844,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 845,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 846,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 847,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 848,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 849,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 850,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 851,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 852,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 853,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 854,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 855,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 856,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 857,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 858,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 859,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 860,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 861,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 862,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 863,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 864,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 865,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 866,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 867,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 868,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 10, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 869,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 870,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 871,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 872,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 873,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 874,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 875,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 876,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 877,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 3, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 878,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 879,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 880,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 881,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 3, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 882,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 883,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 884,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 885,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 886,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 887,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 888,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 889,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 890,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 891,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 892,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 893,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 894,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 895,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 896,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 897,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 898,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 899,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 900,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 8, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 901,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 902,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 903,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 2, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 904,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 905,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 906,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 907,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 908,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 909,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 910,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 911,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 912,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 913,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 914,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 915,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 916,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 1, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 917,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 918,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 919,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 920,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 921,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 922,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 923,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 924,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 925,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 926,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 927,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 928,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 929,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 930,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 931,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 932,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 933,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 934,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 935,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 936,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 937,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 938,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 939,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 940,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 941,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 942,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 943,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 944,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 945,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 946,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 9, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 947,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 948,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 949,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 950,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 951,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 13, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 952,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 953,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 954,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 955,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 956,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 957,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 958,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 959,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 960,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 961,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 962,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 963,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 964,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 965,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 966,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 967,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 968,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 969,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 970,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 971,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 972,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 973,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 974,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 12, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 975,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 976,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 977,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 978,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 979,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 980,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 981,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 982,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 983,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 984,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 985,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 986,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 987,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 988,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 989,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 990,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 991,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 992,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 993,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 994,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 12, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 995,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 9, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 996,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 997,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 998,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 999,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1000,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1001,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1002,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1003,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1004,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1005,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1006,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1007,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1008,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1009,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1010,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 6, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1011,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1012,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1013,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1014,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1015,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1016,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1017,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1018,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1019,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1020,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1021,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1022,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1023,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1024,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1025,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1026,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1027,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1028,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1029,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1030,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1031,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1032,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1033,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1034,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1035,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1036,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1037,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1038,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 11, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1039,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1040,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1041,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 1, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1042,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1043,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1044,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1045,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1046,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1047,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1048,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1049,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1050,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 12, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1051,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1052,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1053,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1054,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1055,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1056,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1057,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1058,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 12, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1059,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1060,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1061,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1062,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1063,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1064,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1065,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1066,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 6, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1067,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1068,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1069,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1070,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1071,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1072,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1073,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1074,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1075,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1076,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1077,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1078,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1079,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1080,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1081,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1082,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1083,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1084,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1085,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1086,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1087,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1088,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1089,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1090,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1091,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 6, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1092,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1093,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 0, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1094,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1095,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1096,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1097,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1098,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1099,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 7, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 8, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 9, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 2, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 14, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 7, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 0, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 0, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 9, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 10, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 5, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 4, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 14, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 6, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 2, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 11, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 3, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 3, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 0, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 6, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 5, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 0, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 6, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 9, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 14, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 9, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 15, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 0, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 2, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 13, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 12, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 12, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 13, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1663,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1664,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1665,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1666,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1667,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1668,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1669,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1670,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1671,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 15, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1672,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1673,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1674,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1675,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1676,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1677,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1678,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1679,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1680,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1681,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1682,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1683,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1684,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1685,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1686,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1687,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1688,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1689,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1690,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1691,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1692,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1693,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1694,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1695,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1696,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 4, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1697,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1698,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1699,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1700,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1701,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1702,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1703,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1704,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1705,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1706,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1707,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1708,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1709,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1710,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1711,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1712,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1713,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1714,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 7, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1715,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1716,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1717,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1718,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1719,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1720,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1721,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 15, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1722,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1723,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1724,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1725,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1726,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1727,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1728,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1729,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 6, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1730,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1731,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1732,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 9, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1733,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1734,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1735,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1736,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1737,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1738,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1739,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1740,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1741,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1742,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1743,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1744,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1745,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1746,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1747,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1748,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1749,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1750,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1751,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1752,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1753,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1754,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1755,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1756,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1757,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1758,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1759,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1760,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 2, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1761,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 7, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1762,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1763,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1764,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1765,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1766,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1767,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1768,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1769,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1770,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1771,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1772,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1773,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1774,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1775,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1776,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1777,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1778,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 8, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1779,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1780,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1781,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1782,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1783,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1784,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1785,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1786,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1787,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1788,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1789,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1790,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1791,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1792,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1793,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1794,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1795,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1796,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1797,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 9, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1798,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1799,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1800,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1801,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1802,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1803,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1804,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1805,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1806,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 11, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1807,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1808,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1809,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1810,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1811,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1812,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1813,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1814,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1815,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1816,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1817,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1818,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1819,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1820,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1821,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1822,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 7, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1823,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1824,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1825,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 4, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1826,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1827,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1828,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1829,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1830,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1831,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1832,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1833,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1834,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1835,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1836,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1837,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1838,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1839,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1840,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 15, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1841,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1842,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1843,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1844,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1845,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1846,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1847,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1848,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1849,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1850,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1851,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1852,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1853,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1854,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1855,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1856,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1857,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1858,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1859,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1860,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1861,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1862,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1863,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1864,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1865,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1866,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1867,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1868,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1869,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1870,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1871,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1872,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1873,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1874,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1875,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1876,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1877,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1878,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1879,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1880,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1881,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1882,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1883,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1884,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 6, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1885,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1886,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1887,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 3, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1888,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1889,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1890,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1891,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1892,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1893,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1894,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1895,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1896,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1897,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1898,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1899,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1900,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1901,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1902,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1903,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1904,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 9, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1905,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1906,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1907,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1908,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1909,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 5, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1910,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1911,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1912,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1913,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1914,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1915,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 5, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1916,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1917,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1918,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 11, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1919,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1920,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1921,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1922,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1923,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1924,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1925,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1926,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1927,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1928,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1929,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1930,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1931,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1932,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1933,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1934,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1935,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1936,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1937,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1938,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1939,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1940,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1941,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1942,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1943,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1944,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1945,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1946,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1947,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 0, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1948,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1949,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1950,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 0, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1951,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1952,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1953,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1954,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1955,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1956,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 2, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1957,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1958,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1959,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1960,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1961,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1962,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1963,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1964,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 14, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1965,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1966,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1967,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1968,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1969,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1970,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1971,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1972,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1973,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1974,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1975,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1976,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1977,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1978,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 1, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1979,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1980,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 13, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1981,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0001; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1982,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1983,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1984,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1985,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1986,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1987,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1988,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1989,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1990,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1991,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1992,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1993,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1994,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1995,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1996,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1997,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1998,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 1999,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2000,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 4, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2001,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2002,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2003,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2004,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2005,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2006,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2007,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2008,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2009,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2010,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2011,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2012,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2013,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2014,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2015,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2016,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2017,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2018,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2019,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2020,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2021,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2022,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2023,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2024,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2025,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2026,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2027,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2028,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 14, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2029,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2030,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2031,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2032,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2033,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2034,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2035,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 1, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2036,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 5, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2037,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2038,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2039,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2040,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 0, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2041,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2042,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2043,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2044,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2045,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2046,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2047,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2048,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2049,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2050,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2051,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2052,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2053,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2054,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2055,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2056,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2057,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2058,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2059,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2060,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2061,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2062,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2063,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2064,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2065,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2066,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2067,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2068,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2069,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2070,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2071,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2072,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2073,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2074,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 1, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2075,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2076,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2077,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2078,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2079,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2080,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2081,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2082,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2083,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2084,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2085,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2086,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2087,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2088,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2089,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2090,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2091,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2092,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2093,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2094,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2095,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 8, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2096,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2097,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2098,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2099,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 8, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 9, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 10, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 3, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 1, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 6, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 13, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 8, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 6, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 9, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 9, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0100; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 15, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 3, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 14, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 3, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 9, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 7, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 3, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 8, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 10, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 1, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 1, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 13, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 15, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 2, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 15, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 14, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 0, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 2, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1100; // Expected: {'sum': 14, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 5, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 0, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 3, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 4, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 4, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 4, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 5, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 0, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2663,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2664,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2665,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 14, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2666,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2667,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2668,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2669,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2670,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2671,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2672,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2673,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2674,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2675,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2676,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2677,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2678,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2679,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2680,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2681,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2682,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2683,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2684,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2685,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2686,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2687,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2688,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2689,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2690,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2691,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2692,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2693,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 4, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2694,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2695,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2696,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2697,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2698,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2699,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 9, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2700,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 8, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2701,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2702,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2703,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2704,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2705,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2706,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2707,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2708,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2709,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2710,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2711,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2712,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2713,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2714,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2715,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2716,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 3, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2717,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2718,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2719,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2720,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2721,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2722,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 12, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2723,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2724,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2725,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2726,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2727,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2728,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2729,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2730,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2731,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2732,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 0, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2733,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2734,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2735,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2736,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2737,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2738,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2739,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2740,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2741,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2742,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2743,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 0, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2744,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2745,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2746,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 14, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2747,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2748,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2749,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2750,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2751,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2752,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2753,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2754,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2755,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2756,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2757,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2758,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2759,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2760,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2761,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2762,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2763,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2764,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2765,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2766,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2767,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2768,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2769,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 2, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2770,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2771,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2772,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2773,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2774,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2775,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2776,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2777,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2778,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2779,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2780,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 4, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2781,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2782,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2783,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2784,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2785,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2786,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2787,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2788,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2789,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2790,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2791,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2792,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2793,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2794,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2795,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2796,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2797,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2798,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2799,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2800,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2801,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2802,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2803,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2804,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 14, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2805,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2806,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 3, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2807,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2808,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2809,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2810,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2811,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2812,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2813,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2814,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2815,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2816,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 11, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2817,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2818,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2819,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1001; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2820,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2821,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2822,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2823,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2824,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2825,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2826,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2827,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2828,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2829,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2830,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2831,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2832,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 0, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2833,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2834,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2835,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2836,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2837,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2838,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2839,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2840,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 13, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2841,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2842,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2843,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2844,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2845,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2846,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2847,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2848,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2849,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2850,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b0111; // Expected: {'sum': 15, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2851,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2852,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 14, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2853,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2854,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2855,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2856,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2857,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2858,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2859,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2860,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2861,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2862,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2863,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2864,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 10, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2865,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2866,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2867,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2868,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2869,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2870,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2871,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2872,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2873,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2874,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2875,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2876,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2877,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2878,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2879,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2880,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1110; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2881,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2882,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2883,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 10, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2884,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2885,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2886,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2887,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2888,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2889,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2890,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2891,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2892,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2893,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 11, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2894,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0011; // Expected: {'sum': 11, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2895,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2896,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2897,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2898,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2899,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2900,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2901,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2902,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2903,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2904,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2905,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2906,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2907,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2908,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2909,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2910,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2911,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2912,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2913,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2914,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2915,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b1111; // Expected: {'sum': 14, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2916,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2917,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2918,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0100; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2919,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2920,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2921,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2922,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2923,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2924,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2925,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2926,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2927,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2928,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2929,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2930,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 12, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2931,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2932,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 7, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2933,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 6, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2934,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2935,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2936,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2937,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0111; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2938,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2939,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2940,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2941,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2942,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0100; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2943,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2944,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2945,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2946,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2947,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2948,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2949,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2950,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2951,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2952,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2953,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2954,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0101; c = 4'b0100; // Expected: {'sum': 15, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2955,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2956,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 5, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2957,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2958,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2959,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2960,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2961,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2962,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2963,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2964,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2965,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2966,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2967,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b0011; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2968,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2969,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2970,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2971,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2972,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2973,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2974,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2975,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2976,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2977,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2978,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2979,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2980,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2981,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2982,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2983,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2984,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2985,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2986,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2987,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1010; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2988,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2989,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2990,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2991,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2992,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2993,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2994,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 8, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2995,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2996,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2997,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2998,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 2999,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3000,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3001,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 4, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3002,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3003,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3004,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3005,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3006,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3007,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3008,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3009,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3010,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3011,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3012,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3013,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3014,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3015,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3016,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3017,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3018,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3019,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3020,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3021,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3022,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3023,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 1, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3024,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3025,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 11, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3026,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3027,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3028,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3029,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3030,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 14, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3031,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3032,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3033,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3034,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3035,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3036,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 6, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3037,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3038,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3039,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3040,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 3, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3041,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3042,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3043,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 8, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3044,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3045,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3046,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3047,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3048,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3049,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0111; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3050,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3051,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3052,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3053,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3054,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3055,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3056,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3057,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 2, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3058,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3059,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3060,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3061,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 14, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3062,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3063,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3064,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 7, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3065,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3066,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3067,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3068,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 3, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3069,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1110; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3070,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3071,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3072,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 15, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3073,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3074,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3075,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3076,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3077,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b1011; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3078,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3079,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3080,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3081,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3082,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b0101; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3083,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3084,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3085,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3086,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 7, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3087,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3088,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3089,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3090,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3091,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3092,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3093,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3094,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 13, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3095,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 11, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3096,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3097,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3098,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3099,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3100,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 15, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3101,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3102,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3103,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3104,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3105,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3106,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3107,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3108,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3109,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0101; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3110,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 5, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3111,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3112,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3113,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3114,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3115,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3116,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0111; // Expected: {'sum': 1, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3117,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3118,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 15, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3119,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3120,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3121,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3122,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3123,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3124,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3125,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3126,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3127,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3128,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3129,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3130,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 5, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3131,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3132,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3133,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3134,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3135,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3136,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3137,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3138,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3139,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0111; c = 4'b1001; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3140,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3141,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3142,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3143,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3144,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3145,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0110; c = 4'b1111; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3146,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3147,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 14, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3148,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 13, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3149,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3150,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b0111; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3151,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3152,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3153,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3154,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3155,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3156,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3157,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3158,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3159,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3160,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b1101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3161,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3162,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3163,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3164,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3165,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3166,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b0010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3167,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3168,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3169,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b0000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3170,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 11, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3171,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3172,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3173,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 13, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3174,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 2, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3175,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3176,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3177,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 15, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3178,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3179,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b0100; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3180,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1001; c = 4'b0010; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3181,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3182,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3183,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 10, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3184,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3185,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3186,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3187,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3188,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 7, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3189,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3190,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3191,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3192,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3193,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3194,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3195,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3196,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3197,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3198,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3199,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 10, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3200,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3201,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3202,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0100; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3203,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3204,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3205,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1111; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3206,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3207,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3208,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3209,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3210,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3211,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 4, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3212,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3213,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3214,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3215,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3216,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3217,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3218,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3219,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3220,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 5, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3221,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 7, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3222,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3223,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3224,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3225,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 2, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3226,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3227,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 14, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3228,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3229,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3230,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3231,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1010; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3232,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3233,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1010; c = 4'b1011; // Expected: {'sum': 9, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3234,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3235,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3236,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3237,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3238,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3239,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3240,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3241,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3242,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b0111; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3243,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3244,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3245,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3246,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3247,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3248,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3249,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3250,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1111; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3251,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3252,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b0001; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3253,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 14, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3254,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3255,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 3, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3256,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3257,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3258,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 9, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3259,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3260,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3261,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3262,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3263,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3264,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3265,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 5, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3266,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1010; c = 4'b0011; // Expected: {'sum': 10, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3267,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b0000; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3268,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3269,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3270,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 12, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3271,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3272,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0111; // Expected: {'sum': 6, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3273,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3274,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3275,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3276,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 15, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3277,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3278,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b1100; // Expected: {'sum': 5, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3279,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 9, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3280,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3281,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3282,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b0001; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3283,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b0000; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3284,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3285,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b0110; // Expected: {'sum': 2, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3286,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 13, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3287,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0110; c = 4'b1101; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3288,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3289,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1000; c = 4'b1100; // Expected: {'sum': 12, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1000; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3290,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3291,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3292,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3293,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3294,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1011; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3295,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3296,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3297,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3298,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3299,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3300,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3301,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0011; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3302,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3303,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b0110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3304,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0111; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3305,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3306,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3307,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3308,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3309,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0011; c = 4'b1101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3310,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3311,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3312,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3313,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 4, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3314,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3315,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b0000; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3316,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3317,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3318,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3319,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3320,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3321,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3322,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3323,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3324,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3325,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1010; c = 4'b0111; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1010; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3326,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3327,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3328,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3329,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 12, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3330,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 3, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3331,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3332,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1011; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3333,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3334,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3335,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3336,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1010; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3337,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3338,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 5, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3339,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0011; c = 4'b0010; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3340,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3341,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3342,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3343,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1100; c = 4'b1010; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1100; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3344,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b0110; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3345,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3346,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3347,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3348,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 4, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3349,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3350,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3351,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 2, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3352,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3353,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 5, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3354,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 9, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3355,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3356,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b0101; // Expected: {'sum': 3, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3357,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3358,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 15, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3359,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3360,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3361,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3362,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3363,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3364,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3365,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1110; c = 4'b1011; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1110; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3366,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3367,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3368,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b1100; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3369,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3370,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 11, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3371,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b1001; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3372,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3373,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1101; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3374,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3375,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3376,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3377,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1111; c = 4'b1000; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3378,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 7, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3379,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0101; c = 4'b1110; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3380,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b1100; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3381,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3382,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 10, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3383,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b1111; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3384,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3385,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 12, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3386,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1000; c = 4'b1001; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3387,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0100; c = 4'b1000; // Expected: {'sum': 0, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0100; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3388,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1000; c = 4'b0100; // Expected: {'sum': 6, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3389,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0011; // Expected: {'sum': 2, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3390,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 10, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3391,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0101; c = 4'b1111; // Expected: {'sum': 9, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3392,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0001; // Expected: {'sum': 1, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3393,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0010; c = 4'b1100; // Expected: {'sum': 12, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0010; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3394,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 6, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3395,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3396,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0000; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0000; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3397,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3398,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1110; c = 4'b1101; // Expected: {'sum': 13, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1110; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3399,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1100; c = 4'b1101; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3400,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3401,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 0, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3402,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 9, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3403,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3404,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3405,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3406,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3407,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3408,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3409,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3410,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3411,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3412,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 8, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3413,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0011; c = 4'b0110; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3414,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3415,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0100; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3416,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0001; // Expected: {'sum': 13, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3417,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1101; // Expected: {'sum': 3, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3418,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3419,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3420,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3421,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3422,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1100; c = 4'b0011; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1100; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3423,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3424,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3425,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0000; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0000; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3426,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0110; c = 4'b1001; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3427,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3428,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b0100; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3429,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1111; c = 4'b0001; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3430,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3431,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0001; c = 4'b1000; // Expected: {'sum': 1, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3432,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3433,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0011; c = 4'b0001; // Expected: {'sum': 11, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0011; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3434,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3435,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3436,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0001; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3437,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3438,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 7, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3439,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 5, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3440,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0011; // Expected: {'sum': 0, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3441,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1011; c = 4'b1010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3442,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0001; c = 4'b0000; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3443,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0000; c = 4'b1111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0000; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3444,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0111; // Expected: {'sum': 5, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3445,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3446,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3447,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3448,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 3, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3449,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3450,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3451,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3452,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3453,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b0001; // Expected: {'sum': 2, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3454,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3455,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1001; // Expected: {'sum': 0, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3456,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3457,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 4, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3458,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3459,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0110; c = 4'b0101; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3460,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3461,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3462,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3463,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3464,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1110; c = 4'b0000; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3465,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0011; c = 4'b1011; // Expected: {'sum': 11, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0011; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3466,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3467,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1111; c = 4'b0110; // Expected: {'sum': 15, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1111; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3468,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0101; c = 4'b0011; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3469,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3470,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b0100; // Expected: {'sum': 1, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3471,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1111; c = 4'b1011; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3472,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1001; c = 4'b1101; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3473,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0011; c = 4'b1110; // Expected: {'sum': 7, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3474,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3475,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0100; c = 4'b1011; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3476,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3477,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b0001; // Expected: {'sum': 13, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3478,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 12, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3479,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 12, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3480,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 5, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3481,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 4, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3482,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1111; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3483,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3484,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b1001; // Expected: {'sum': 1, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3485,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 0, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3486,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 3, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3487,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3488,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3489,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3490,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3491,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b1100; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3492,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3493,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1110; // Expected: {'sum': 7, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3494,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 14, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3495,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0111; c = 4'b1011; // Expected: {'sum': 15, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0111; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3496,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3497,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 7, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3498,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3499,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b0000; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3500,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 13, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3501,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b0000; // Expected: {'sum': 4, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3502,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b1100; // Expected: {'sum': 13, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3503,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1011; c = 4'b1110; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1011; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3504,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 4, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3505,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3506,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3507,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b1100; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3508,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3509,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3510,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3511,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3512,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0110; // Expected: {'sum': 6, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3513,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3514,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0011; // Expected: {'sum': 9, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3515,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1100; c = 4'b0110; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3516,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0001; c = 4'b1010; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3517,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1101; c = 4'b0011; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1101; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3518,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0111; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3519,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3520,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3521,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3522,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3523,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3524,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b0100; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3525,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3526,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0011; c = 4'b0100; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0011; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3527,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 5, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3528,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 11, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3529,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1010; c = 4'b1010; // Expected: {'sum': 6, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3530,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 10, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3531,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1011; c = 4'b0010; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1011; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3532,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 4, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3533,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3534,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0000; c = 4'b0101; // Expected: {'sum': 9, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3535,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0111; c = 4'b0000; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0111; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3536,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0111; c = 4'b0011; // Expected: {'sum': 6, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0111; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3537,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b1010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3538,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1001; c = 4'b0101; // Expected: {'sum': 11, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1001; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3539,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1111; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3540,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1010; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1010; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3541,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b0101; // Expected: {'sum': 2, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3542,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0010; c = 4'b1011; // Expected: {'sum': 8, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0010; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3543,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0101; c = 4'b1100; // Expected: {'sum': 6, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0101; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3544,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b0010; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3545,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1110; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1110; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3546,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 12, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3547,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3548,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3549,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0110; c = 4'b1100; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0110; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3550,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1101; c = 4'b0100; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1101; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3551,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0001; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3552,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 8, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3553,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0110; c = 4'b0010; // Expected: {'sum': 2, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0110; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3554,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b1110; // Expected: {'sum': 4, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3555,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0100; c = 4'b1111; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0100; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3556,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1001; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3557,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0010; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3558,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1111; // Expected: {'sum': 9, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3559,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1111; c = 4'b1100; // Expected: {'sum': 15, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3560,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1101; c = 4'b0101; // Expected: {'sum': 5, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1101; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3561,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0011; c = 4'b1010; // Expected: {'sum': 6, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0011; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3562,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1101; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3563,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b1110; c = 4'b1000; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b1110; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3564,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3565,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1000; // Expected: {'sum': 12, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3566,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0101; c = 4'b1010; // Expected: {'sum': 11, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0101; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3567,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1001; c = 4'b0000; // Expected: {'sum': 8, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1001; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3568,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0100; c = 4'b1001; // Expected: {'sum': 0, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0100; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3569,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0111; c = 4'b1100; // Expected: {'sum': 5, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0111; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3570,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0111; c = 4'b1000; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0111; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3571,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0111; c = 4'b1010; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0111; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3572,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b0001; // Expected: {'sum': 5, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3573,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1100; c = 4'b1011; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1100; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3574,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1100; c = 4'b0010; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3575,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 8, 'carry': 7}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3576,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b0001; c = 4'b1111; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b0001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3577,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0010; c = 4'b0000; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0010; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3578,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1111; c = 4'b1001; // Expected: {'sum': 13, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1111; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3579,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0001; c = 4'b1001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0001; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3580,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1110; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3581,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1101; c = 4'b1101; // Expected: {'sum': 9, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1101; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3582,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0011; b = 4'b0001; c = 4'b1101; // Expected: {'sum': 15, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0011; b = 4'b0001; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3583,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3584,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1111; c = 4'b1110; // Expected: {'sum': 4, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1111; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3585,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 4, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 2, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3586,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1100; c = 4'b0000; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1100; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3587,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3588,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3589,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 10, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3590,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1110; c = 4'b0101; // Expected: {'sum': 1, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1110; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3591,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1001; c = 4'b1011; // Expected: {'sum': 8, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1001; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3592,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3593,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 11, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3594,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3595,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0100; c = 4'b0100; // Expected: {'sum': 6, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0100; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3596,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1110; c = 4'b0011; // Expected: {'sum': 2, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1110; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3597,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 3, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3598,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1000; c = 4'b0101; // Expected: {'sum': 6, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1000; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3599,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b0010; c = 4'b0001; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b0010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3600,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b0110; // Expected: {'sum': 10, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3601,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0001; c = 4'b1110; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3602,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1010; // Expected: {'sum': 0, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3603,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1011; c = 4'b0111; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1011; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3604,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3605,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b0110; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3606,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 11, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3607,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b1001; // Expected: {'sum': 9, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3608,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 1, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3609,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b1001; c = 4'b1110; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b1001; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3610,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1011; c = 4'b0000; // Expected: {'sum': 13, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3611,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3612,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0100; c = 4'b0110; // Expected: {'sum': 8, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0100; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3613,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b1111; c = 4'b1111; // Expected: {'sum': 10, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b1111; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3614,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3615,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1000; c = 4'b1101; // Expected: {'sum': 3, 'carry': 12}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1000; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3616,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3617,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1101; b = 4'b1001; c = 4'b1100; // Expected: {'sum': 8, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1101; b = 4'b1001; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3618,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1111; c = 4'b1101; // Expected: {'sum': 10, 'carry': 13}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3619,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 14, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3620,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1001; b = 4'b0010; c = 4'b1000; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1001; b = 4'b0010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3621,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1100; c = 4'b0001; // Expected: {'sum': 12, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1100; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3622,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0111; c = 4'b0101; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0111; c = 4'b0101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3623,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b1000; c = 4'b0110; // Expected: {'sum': 10, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b1000; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3624,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3625,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0101; c = 4'b0110; // Expected: {'sum': 6, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3626,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1101; c = 4'b1011; // Expected: {'sum': 14, 'carry': 9}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1101; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3627,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1000; // Expected: {'sum': 12, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3628,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0000; c = 4'b0111; // Expected: {'sum': 6, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3629,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 6, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0000; c = 4'b0010; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0000; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3630,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1100; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3631,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0111; c = 4'b1101; // Expected: {'sum': 1, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0111; c = 4'b1101; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3632,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b0110; c = 4'b0000; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b0110; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3633,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1010; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 10, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1010; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3634,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b1010; c = 4'b1001; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b1010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3635,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1011; c = 4'b1000; // Expected: {'sum': 1, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1011; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3636,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0101; c = 4'b0111; // Expected: {'sum': 10, 'carry': 5}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0101; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3637,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 10, 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0000; b = 4'b0101; c = 4'b0010; // Expected: {'sum': 7, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0000; b = 4'b0101; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3638,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0100; c = 4'b0010; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0100; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3639,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1100; b = 4'b1010; c = 4'b1000; // Expected: {'sum': 14, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1100; b = 4'b1010; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3640,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0101; b = 4'b0110; c = 4'b1110; // Expected: {'sum': 13, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0101; b = 4'b0110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3641,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 13, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 5, 'carry': 10}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3642,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 5, 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0001; b = 4'b1000; c = 4'b0111; // Expected: {'sum': 14, 'carry': 1}
        #10;
        $display("Test %0d: Inputs: a = 4'b0001; b = 4'b1000; c = 4'b0111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3643,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 14, 
                 
                 1
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b0001; c = 4'b0010; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b0001; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3644,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b1001; c = 4'b1111; // Expected: {'sum': 0, 'carry': 15}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b1001; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3645,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 0, 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b0110; // Expected: {'sum': 9, 'carry': 6}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3646,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 9, 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b1001; // Expected: {'sum': 3, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3647,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 3, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1110; b = 4'b1000; c = 4'b1110; // Expected: {'sum': 8, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b1110; b = 4'b1000; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3648,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b0001; c = 4'b0110; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b0001; c = 4'b0110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3649,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b0011; c = 4'b0000; // Expected: {'sum': 1, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b0011; c = 4'b0000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3650,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 1, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0100; b = 4'b0000; c = 4'b1011; // Expected: {'sum': 15, 'carry': 0}
        #10;
        $display("Test %0d: Inputs: a = 4'b0100; b = 4'b0000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3651,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1110; c = 4'b1110; // Expected: {'sum': 7, 'carry': 14}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1110; c = 4'b1110; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3652,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1011; b = 4'b1011; c = 4'b1111; // Expected: {'sum': 15, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1011; b = 4'b1011; c = 4'b1111; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3653,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0010; b = 4'b1101; c = 4'b1000; // Expected: {'sum': 7, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b0010; b = 4'b1101; c = 4'b1000; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3654,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 7, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0001; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3655,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1000; c = 4'b0011; // Expected: {'sum': 12, 'carry': 3}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1000; c = 4'b0011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3656,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b0010; c = 4'b0010; // Expected: {'sum': 8, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b0010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3657,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 8, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0111; b = 4'b1010; c = 4'b0010; // Expected: {'sum': 15, 'carry': 2}
        #10;
        $display("Test %0d: Inputs: a = 4'b0111; b = 4'b1010; c = 4'b0010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3658,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1110; c = 4'b1001; // Expected: {'sum': 15, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1110; c = 4'b1001; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3659,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 15, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b0110; b = 4'b0000; c = 4'b0100; // Expected: {'sum': 2, 'carry': 4}
        #10;
        $display("Test %0d: Inputs: a = 4'b0110; b = 4'b0000; c = 4'b0100; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3660,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 2, 
                 
                 4
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1111; b = 4'b1000; c = 4'b1011; // Expected: {'sum': 12, 'carry': 11}
        #10;
        $display("Test %0d: Inputs: a = 4'b1111; b = 4'b1000; c = 4'b1011; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3661,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 12, 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 4'b1000; b = 4'b1001; c = 4'b1010; // Expected: {'sum': 11, 'carry': 8}
        #10;
        $display("Test %0d: Inputs: a = 4'b1000; b = 4'b1001; c = 4'b1010; | Outputs: sum=%b, carry=%b | Expected: sum=%d, carry=%d",
                 3662,
                 
                 sum, 
                 
                 carry
                 , 
                 
                 11, 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule