
`timescale 1ns / 1ps

module tb_N6_array_multiplier;

    // Parameters
    
    parameter N = 6;
    
     
    // Inputs
    
    reg  [5:0] A;
    
    reg  [5:0] B;
    
    
    // Outputs
    
    wire   P;
    
    
    // Instantiate the Unit Under Test (UUT)
    array_multiplier  #( N ) uut (
        
        .A(A),
        
        .B(B),
        
        
        .P(P)
        
    );

    // Clock generation 
    

    
    
    initial begin
        // Initialize Inputs
        
        A = 0;
        
        B = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 A = 6'b011111; B = 6'b101011; // Expected: {'P': 1333}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 0,
                 
                 P
                 , 
                 
                 1333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b011001; // Expected: {'P': 425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1,
                 
                 P
                 , 
                 
                 425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b001111; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000001; // Expected: {'P': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 3,
                 
                 P
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111100; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 4,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b011001; // Expected: {'P': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 5,
                 
                 P
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001110; // Expected: {'P': 476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 6,
                 
                 P
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b111110; // Expected: {'P': 2108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 7,
                 
                 P
                 , 
                 
                 2108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b110010; // Expected: {'P': 2300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 8,
                 
                 P
                 , 
                 
                 2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100010; // Expected: {'P': 1428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 9,
                 
                 P
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b111101; // Expected: {'P': 244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 10,
                 
                 P
                 , 
                 
                 244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b000101; // Expected: {'P': 290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 11,
                 
                 P
                 , 
                 
                 290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 12,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b001110; // Expected: {'P': 812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 13,
                 
                 P
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b100011; // Expected: {'P': 1995}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 14,
                 
                 P
                 , 
                 
                 1995
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b001000; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 15,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b011000; // Expected: {'P': 864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 16,
                 
                 P
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b111000; // Expected: {'P': 952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 17,
                 
                 P
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001111; // Expected: {'P': 510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 18,
                 
                 P
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b111001; // Expected: {'P': 3249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 19,
                 
                 P
                 , 
                 
                 3249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b111010; // Expected: {'P': 2088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 20,
                 
                 P
                 , 
                 
                 2088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b001010; // Expected: {'P': 620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 21,
                 
                 P
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110100; // Expected: {'P': 2028}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 22,
                 
                 P
                 , 
                 
                 2028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001100; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 23,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b000011; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 24,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b010110; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 25,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b001111; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 26,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100101; // Expected: {'P': 481}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 27,
                 
                 P
                 , 
                 
                 481
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011100; // Expected: {'P': 1764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 28,
                 
                 P
                 , 
                 
                 1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110000; // Expected: {'P': 1536}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 29,
                 
                 P
                 , 
                 
                 1536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b011110; // Expected: {'P': 870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 30,
                 
                 P
                 , 
                 
                 870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b010111; // Expected: {'P': 414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 31,
                 
                 P
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b101010; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 32,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b011110; // Expected: {'P': 1740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 33,
                 
                 P
                 , 
                 
                 1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b100101; // Expected: {'P': 1332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 34,
                 
                 P
                 , 
                 
                 1332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000111; // Expected: {'P': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 35,
                 
                 P
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b010001; // Expected: {'P': 935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 36,
                 
                 P
                 , 
                 
                 935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b111111; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 37,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b010100; // Expected: {'P': 1060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 38,
                 
                 P
                 , 
                 
                 1060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011001; // Expected: {'P': 475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 39,
                 
                 P
                 , 
                 
                 475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b011100; // Expected: {'P': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 40,
                 
                 P
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100010; // Expected: {'P': 1258}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 41,
                 
                 P
                 , 
                 
                 1258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b011101; // Expected: {'P': 1305}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 42,
                 
                 P
                 , 
                 
                 1305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 43,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b101011; // Expected: {'P': 1720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 44,
                 
                 P
                 , 
                 
                 1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b010011; // Expected: {'P': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 45,
                 
                 P
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011110; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 46,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b011101; // Expected: {'P': 1682}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 47,
                 
                 P
                 , 
                 
                 1682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b001010; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 48,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b111111; // Expected: {'P': 1071}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 49,
                 
                 P
                 , 
                 
                 1071
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b000100; // Expected: {'P': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 50,
                 
                 P
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b101111; // Expected: {'P': 1410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 51,
                 
                 P
                 , 
                 
                 1410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b010101; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 52,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b001111; // Expected: {'P': 825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 53,
                 
                 P
                 , 
                 
                 825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b011011; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 54,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b000100; // Expected: {'P': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 55,
                 
                 P
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b110011; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 56,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b110010; // Expected: {'P': 2000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 57,
                 
                 P
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b110111; // Expected: {'P': 605}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 58,
                 
                 P
                 , 
                 
                 605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100100; // Expected: {'P': 1476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 59,
                 
                 P
                 , 
                 
                 1476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b011101; // Expected: {'P': 754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 60,
                 
                 P
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b010011; // Expected: {'P': 171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 61,
                 
                 P
                 , 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000100; // Expected: {'P': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 62,
                 
                 P
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b011110; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 63,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b000001; // Expected: {'P': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 64,
                 
                 P
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b001110; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 65,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b111110; // Expected: {'P': 1984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 66,
                 
                 P
                 , 
                 
                 1984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b000001; // Expected: {'P': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 67,
                 
                 P
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b110010; // Expected: {'P': 800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 68,
                 
                 P
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001110; // Expected: {'P': 854}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 69,
                 
                 P
                 , 
                 
                 854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b010110; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 70,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101110; // Expected: {'P': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 71,
                 
                 P
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b001110; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 72,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b110010; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 73,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b000101; // Expected: {'P': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 74,
                 
                 P
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b101101; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 75,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b010010; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 76,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b110100; // Expected: {'P': 676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 77,
                 
                 P
                 , 
                 
                 676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b011100; // Expected: {'P': 868}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 78,
                 
                 P
                 , 
                 
                 868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000100; // Expected: {'P': 152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 79,
                 
                 P
                 , 
                 
                 152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000001; // Expected: {'P': 3}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 80,
                 
                 P
                 , 
                 
                 3
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b010110; // Expected: {'P': 836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 81,
                 
                 P
                 , 
                 
                 836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b100100; // Expected: {'P': 1908}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 82,
                 
                 P
                 , 
                 
                 1908
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b101010; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 83,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101001; // Expected: {'P': 1435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 84,
                 
                 P
                 , 
                 
                 1435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b101000; // Expected: {'P': 2480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 85,
                 
                 P
                 , 
                 
                 2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b010001; // Expected: {'P': 357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 86,
                 
                 P
                 , 
                 
                 357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b001100; // Expected: {'P': 348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 87,
                 
                 P
                 , 
                 
                 348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 88,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b110011; // Expected: {'P': 2091}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 89,
                 
                 P
                 , 
                 
                 2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b111100; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 90,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010100; // Expected: {'P': 620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 91,
                 
                 P
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b001010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 92,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b010010; // Expected: {'P': 612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 93,
                 
                 P
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000100; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 94,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b101010; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 95,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b000010; // Expected: {'P': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 96,
                 
                 P
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b001100; // Expected: {'P': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 97,
                 
                 P
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b010000; // Expected: {'P': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 98,
                 
                 P
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b101100; // Expected: {'P': 1276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 99,
                 
                 P
                 , 
                 
                 1276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100100; // Expected: {'P': 972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 100,
                 
                 P
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b100110; // Expected: {'P': 1216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 101,
                 
                 P
                 , 
                 
                 1216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b010000; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 102,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b111111; // Expected: {'P': 2835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 103,
                 
                 P
                 , 
                 
                 2835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b011001; // Expected: {'P': 1250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 104,
                 
                 P
                 , 
                 
                 1250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b111110; // Expected: {'P': 3658}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 105,
                 
                 P
                 , 
                 
                 3658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b100011; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 106,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b100010; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 107,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b001100; // Expected: {'P': 696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 108,
                 
                 P
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b010010; // Expected: {'P': 810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 109,
                 
                 P
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b100101; // Expected: {'P': 2257}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 110,
                 
                 P
                 , 
                 
                 2257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b110001; // Expected: {'P': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 111,
                 
                 P
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b010111; // Expected: {'P': 1265}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 112,
                 
                 P
                 , 
                 
                 1265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b000101; // Expected: {'P': 95}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 113,
                 
                 P
                 , 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b000100; // Expected: {'P': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 114,
                 
                 P
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b010110; // Expected: {'P': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 115,
                 
                 P
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b111001; // Expected: {'P': 2223}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 116,
                 
                 P
                 , 
                 
                 2223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b100111; // Expected: {'P': 2379}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 117,
                 
                 P
                 , 
                 
                 2379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b100111; // Expected: {'P': 1014}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 118,
                 
                 P
                 , 
                 
                 1014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b011100; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 119,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b010111; // Expected: {'P': 483}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 120,
                 
                 P
                 , 
                 
                 483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001100; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 121,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b001011; // Expected: {'P': 143}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 122,
                 
                 P
                 , 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b100001; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 123,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b000010; // Expected: {'P': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 124,
                 
                 P
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b101101; // Expected: {'P': 1710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 125,
                 
                 P
                 , 
                 
                 1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b101011; // Expected: {'P': 1290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 126,
                 
                 P
                 , 
                 
                 1290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100101; // Expected: {'P': 1702}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 127,
                 
                 P
                 , 
                 
                 1702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b110001; // Expected: {'P': 1225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 128,
                 
                 P
                 , 
                 
                 1225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b101101; // Expected: {'P': 2745}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 129,
                 
                 P
                 , 
                 
                 2745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b000110; // Expected: {'P': 348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 130,
                 
                 P
                 , 
                 
                 348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b010001; // Expected: {'P': 765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 131,
                 
                 P
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000001; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 132,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b010100; // Expected: {'P': 1140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 133,
                 
                 P
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b101000; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 134,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b110110; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 135,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 136,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000010; // Expected: {'P': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 137,
                 
                 P
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b010101; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 138,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111101; // Expected: {'P': 2806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 139,
                 
                 P
                 , 
                 
                 2806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b100100; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 140,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001010; // Expected: {'P': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 141,
                 
                 P
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100001; // Expected: {'P': 627}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 142,
                 
                 P
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010010; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 143,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100010; // Expected: {'P': 646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 144,
                 
                 P
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111011; // Expected: {'P': 944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 145,
                 
                 P
                 , 
                 
                 944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b010010; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 146,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 147,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b100100; // Expected: {'P': 1044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 148,
                 
                 P
                 , 
                 
                 1044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b011010; // Expected: {'P': 1430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 149,
                 
                 P
                 , 
                 
                 1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b001000; // Expected: {'P': 392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 150,
                 
                 P
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b001111; // Expected: {'P': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 151,
                 
                 P
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b000100; // Expected: {'P': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 152,
                 
                 P
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b000010; // Expected: {'P': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 153,
                 
                 P
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b111100; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 154,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b001000; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 155,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b010001; // Expected: {'P': 323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 156,
                 
                 P
                 , 
                 
                 323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b010000; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 157,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010110; // Expected: {'P': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 158,
                 
                 P
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b111011; // Expected: {'P': 1416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 159,
                 
                 P
                 , 
                 
                 1416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b111011; // Expected: {'P': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 160,
                 
                 P
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b010100; // Expected: {'P': 580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 161,
                 
                 P
                 , 
                 
                 580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011000; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 162,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b001110; // Expected: {'P': 266}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 163,
                 
                 P
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b010001; // Expected: {'P': 612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 164,
                 
                 P
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b011011; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 165,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b011011; // Expected: {'P': 351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 166,
                 
                 P
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b111101; // Expected: {'P': 2013}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 167,
                 
                 P
                 , 
                 
                 2013
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000011; // Expected: {'P': 105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 168,
                 
                 P
                 , 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010010; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 169,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b001100; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 170,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b111111; // Expected: {'P': 3276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 171,
                 
                 P
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b000001; // Expected: {'P': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 172,
                 
                 P
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b111001; // Expected: {'P': 1710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 173,
                 
                 P
                 , 
                 
                 1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b110011; // Expected: {'P': 1479}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 174,
                 
                 P
                 , 
                 
                 1479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b111111; // Expected: {'P': 441}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 175,
                 
                 P
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111011; // Expected: {'P': 2714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 176,
                 
                 P
                 , 
                 
                 2714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b101001; // Expected: {'P': 1271}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 177,
                 
                 P
                 , 
                 
                 1271
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b101100; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 178,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b010100; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 179,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b011101; // Expected: {'P': 1595}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 180,
                 
                 P
                 , 
                 
                 1595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b111100; // Expected: {'P': 1560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 181,
                 
                 P
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b010000; // Expected: {'P': 784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 182,
                 
                 P
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 183,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b101011; // Expected: {'P': 1892}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 184,
                 
                 P
                 , 
                 
                 1892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b001010; // Expected: {'P': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 185,
                 
                 P
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b111001; // Expected: {'P': 2109}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 186,
                 
                 P
                 , 
                 
                 2109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b001010; // Expected: {'P': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 187,
                 
                 P
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b111000; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 188,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001101; // Expected: {'P': 299}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 189,
                 
                 P
                 , 
                 
                 299
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b011110; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 190,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101101; // Expected: {'P': 2205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 191,
                 
                 P
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b101111; // Expected: {'P': 1786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 192,
                 
                 P
                 , 
                 
                 1786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b010111; // Expected: {'P': 736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 193,
                 
                 P
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b011101; // Expected: {'P': 1276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 194,
                 
                 P
                 , 
                 
                 1276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b011100; // Expected: {'P': 952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 195,
                 
                 P
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b110111; // Expected: {'P': 2310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 196,
                 
                 P
                 , 
                 
                 2310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100110; // Expected: {'P': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 197,
                 
                 P
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b000110; // Expected: {'P': 138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 198,
                 
                 P
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010000; // Expected: {'P': 704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 199,
                 
                 P
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000101; // Expected: {'P': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 200,
                 
                 P
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 201,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b110010; // Expected: {'P': 1250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 202,
                 
                 P
                 , 
                 
                 1250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011110; // Expected: {'P': 1530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 203,
                 
                 P
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101110; // Expected: {'P': 2254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 204,
                 
                 P
                 , 
                 
                 2254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110101; // Expected: {'P': 530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 205,
                 
                 P
                 , 
                 
                 530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b011000; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 206,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b110110; // Expected: {'P': 3132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 207,
                 
                 P
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b011011; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 208,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b110100; // Expected: {'P': 1196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 209,
                 
                 P
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b000010; // Expected: {'P': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 210,
                 
                 P
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b011100; // Expected: {'P': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 211,
                 
                 P
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110001; // Expected: {'P': 2744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 212,
                 
                 P
                 , 
                 
                 2744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b011111; // Expected: {'P': 930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 213,
                 
                 P
                 , 
                 
                 930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b101011; // Expected: {'P': 2537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 214,
                 
                 P
                 , 
                 
                 2537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b001101; // Expected: {'P': 572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 215,
                 
                 P
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b100010; // Expected: {'P': 1292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 216,
                 
                 P
                 , 
                 
                 1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100100; // Expected: {'P': 1332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 217,
                 
                 P
                 , 
                 
                 1332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b111110; // Expected: {'P': 2914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 218,
                 
                 P
                 , 
                 
                 2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110001; // Expected: {'P': 1911}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 219,
                 
                 P
                 , 
                 
                 1911
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b010100; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 220,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110110; // Expected: {'P': 1728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 221,
                 
                 P
                 , 
                 
                 1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b110011; // Expected: {'P': 1173}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 222,
                 
                 P
                 , 
                 
                 1173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100000; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 223,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b011001; // Expected: {'P': 275}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 224,
                 
                 P
                 , 
                 
                 275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111010; // Expected: {'P': 522}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 225,
                 
                 P
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b111111; // Expected: {'P': 2142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 226,
                 
                 P
                 , 
                 
                 2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 227,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b111110; // Expected: {'P': 2542}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 228,
                 
                 P
                 , 
                 
                 2542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b101001; // Expected: {'P': 820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 229,
                 
                 P
                 , 
                 
                 820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b010101; // Expected: {'P': 819}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 230,
                 
                 P
                 , 
                 
                 819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110001; // Expected: {'P': 147}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 231,
                 
                 P
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b111011; // Expected: {'P': 1829}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 232,
                 
                 P
                 , 
                 
                 1829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b011010; // Expected: {'P': 1014}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 233,
                 
                 P
                 , 
                 
                 1014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b101100; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 234,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001100; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 235,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b100111; // Expected: {'P': 1326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 236,
                 
                 P
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b110110; // Expected: {'P': 2376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 237,
                 
                 P
                 , 
                 
                 2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b111010; // Expected: {'P': 406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 238,
                 
                 P
                 , 
                 
                 406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b100111; // Expected: {'P': 897}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 239,
                 
                 P
                 , 
                 
                 897
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b011111; // Expected: {'P': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 240,
                 
                 P
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b110101; // Expected: {'P': 2279}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 241,
                 
                 P
                 , 
                 
                 2279
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b111101; // Expected: {'P': 488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 242,
                 
                 P
                 , 
                 
                 488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b101101; // Expected: {'P': 1485}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 243,
                 
                 P
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000110; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 244,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110011; // Expected: {'P': 1530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 245,
                 
                 P
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b100011; // Expected: {'P': 1085}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 246,
                 
                 P
                 , 
                 
                 1085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b001100; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 247,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b001000; // Expected: {'P': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 248,
                 
                 P
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010011; // Expected: {'P': 589}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 249,
                 
                 P
                 , 
                 
                 589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b011101; // Expected: {'P': 1653}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 250,
                 
                 P
                 , 
                 
                 1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b011010; // Expected: {'P': 286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 251,
                 
                 P
                 , 
                 
                 286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b110111; // Expected: {'P': 1155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 252,
                 
                 P
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b010011; // Expected: {'P': 988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 253,
                 
                 P
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b100111; // Expected: {'P': 1482}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 254,
                 
                 P
                 , 
                 
                 1482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111001; // Expected: {'P': 3420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 255,
                 
                 P
                 , 
                 
                 3420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b100010; // Expected: {'P': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 256,
                 
                 P
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b101000; // Expected: {'P': 2160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 257,
                 
                 P
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b110001; // Expected: {'P': 2989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 258,
                 
                 P
                 , 
                 
                 2989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b111110; // Expected: {'P': 1178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 259,
                 
                 P
                 , 
                 
                 1178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b011111; // Expected: {'P': 1271}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 260,
                 
                 P
                 , 
                 
                 1271
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b100101; // Expected: {'P': 1998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 261,
                 
                 P
                 , 
                 
                 1998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b110000; // Expected: {'P': 1968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 262,
                 
                 P
                 , 
                 
                 1968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b000110; // Expected: {'P': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 263,
                 
                 P
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b110010; // Expected: {'P': 1300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 264,
                 
                 P
                 , 
                 
                 1300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b101011; // Expected: {'P': 946}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 265,
                 
                 P
                 , 
                 
                 946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b111101; // Expected: {'P': 1525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 266,
                 
                 P
                 , 
                 
                 1525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b100101; // Expected: {'P': 1591}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 267,
                 
                 P
                 , 
                 
                 1591
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011100; // Expected: {'P': 1428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 268,
                 
                 P
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b011011; // Expected: {'P': 459}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 269,
                 
                 P
                 , 
                 
                 459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b101110; // Expected: {'P': 414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 270,
                 
                 P
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b101100; // Expected: {'P': 572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 271,
                 
                 P
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101001; // Expected: {'P': 656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 272,
                 
                 P
                 , 
                 
                 656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b000010; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 273,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b000010; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 274,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b010011; // Expected: {'P': 741}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 275,
                 
                 P
                 , 
                 
                 741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011000; // Expected: {'P': 456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 276,
                 
                 P
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b010010; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 277,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111000; // Expected: {'P': 2352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 278,
                 
                 P
                 , 
                 
                 2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111111; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 279,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b111100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 280,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b110100; // Expected: {'P': 1924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 281,
                 
                 P
                 , 
                 
                 1924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b110111; // Expected: {'P': 770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 282,
                 
                 P
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b111111; // Expected: {'P': 1953}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 283,
                 
                 P
                 , 
                 
                 1953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b011011; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 284,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b001100; // Expected: {'P': 744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 285,
                 
                 P
                 , 
                 
                 744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b101000; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 286,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 287,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b110100; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 288,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b100010; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 289,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b010001; // Expected: {'P': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 290,
                 
                 P
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b001101; // Expected: {'P': 377}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 291,
                 
                 P
                 , 
                 
                 377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b111001; // Expected: {'P': 2736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 292,
                 
                 P
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000011; // Expected: {'P': 87}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 293,
                 
                 P
                 , 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b110010; // Expected: {'P': 2150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 294,
                 
                 P
                 , 
                 
                 2150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b101101; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 295,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b000100; // Expected: {'P': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 296,
                 
                 P
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b111111; // Expected: {'P': 3213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 297,
                 
                 P
                 , 
                 
                 3213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100111; // Expected: {'P': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 298,
                 
                 P
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b000100; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 299,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b110010; // Expected: {'P': 2050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 300,
                 
                 P
                 , 
                 
                 2050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b010111; // Expected: {'P': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 301,
                 
                 P
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100010; // Expected: {'P': 510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 302,
                 
                 P
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b001011; // Expected: {'P': 682}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 303,
                 
                 P
                 , 
                 
                 682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b101000; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 304,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b001011; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 305,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000101; // Expected: {'P': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 306,
                 
                 P
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b000001; // Expected: {'P': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 307,
                 
                 P
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b001011; // Expected: {'P': 649}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 308,
                 
                 P
                 , 
                 
                 649
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b101100; // Expected: {'P': 1892}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 309,
                 
                 P
                 , 
                 
                 1892
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b001001; // Expected: {'P': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 310,
                 
                 P
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b111100; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 311,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b011011; // Expected: {'P': 675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 312,
                 
                 P
                 , 
                 
                 675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b001010; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 313,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b100011; // Expected: {'P': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 314,
                 
                 P
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b010011; // Expected: {'P': 1102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 315,
                 
                 P
                 , 
                 
                 1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001111; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 316,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b111000; // Expected: {'P': 616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 317,
                 
                 P
                 , 
                 
                 616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b001101; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 318,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b100001; // Expected: {'P': 957}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 319,
                 
                 P
                 , 
                 
                 957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b110000; // Expected: {'P': 2928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 320,
                 
                 P
                 , 
                 
                 2928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b010111; // Expected: {'P': 1449}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 321,
                 
                 P
                 , 
                 
                 1449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111010; // Expected: {'P': 3480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 322,
                 
                 P
                 , 
                 
                 3480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011001; // Expected: {'P': 1175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 323,
                 
                 P
                 , 
                 
                 1175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b000101; // Expected: {'P': 155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 324,
                 
                 P
                 , 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000110; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 325,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011111; // Expected: {'P': 589}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 326,
                 
                 P
                 , 
                 
                 589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b001110; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 327,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101010; // Expected: {'P': 1470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 328,
                 
                 P
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010100; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 329,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b100001; // Expected: {'P': 1617}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 330,
                 
                 P
                 , 
                 
                 1617
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001011; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 331,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b011000; // Expected: {'P': 552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 332,
                 
                 P
                 , 
                 
                 552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101111; // Expected: {'P': 1645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 333,
                 
                 P
                 , 
                 
                 1645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b010001; // Expected: {'P': 340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 334,
                 
                 P
                 , 
                 
                 340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b011000; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 335,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b111101; // Expected: {'P': 2440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 336,
                 
                 P
                 , 
                 
                 2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b001100; // Expected: {'P': 420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 337,
                 
                 P
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b011111; // Expected: {'P': 961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 338,
                 
                 P
                 , 
                 
                 961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b000110; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 339,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b101110; // Expected: {'P': 1426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 340,
                 
                 P
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b100101; // Expected: {'P': 1221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 341,
                 
                 P
                 , 
                 
                 1221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011101; // Expected: {'P': 1827}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 342,
                 
                 P
                 , 
                 
                 1827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b100001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 343,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b110001; // Expected: {'P': 343}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 344,
                 
                 P
                 , 
                 
                 343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b100110; // Expected: {'P': 646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 345,
                 
                 P
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b001111; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 346,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111000; // Expected: {'P': 2576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 347,
                 
                 P
                 , 
                 
                 2576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b101101; // Expected: {'P': 1935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 348,
                 
                 P
                 , 
                 
                 1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b000110; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 349,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b110110; // Expected: {'P': 3186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 350,
                 
                 P
                 , 
                 
                 3186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b111100; // Expected: {'P': 2820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 351,
                 
                 P
                 , 
                 
                 2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b110011; // Expected: {'P': 765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 352,
                 
                 P
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 353,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b101111; // Expected: {'P': 705}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 354,
                 
                 P
                 , 
                 
                 705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100001; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 355,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101001; // Expected: {'P': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 356,
                 
                 P
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b101000; // Expected: {'P': 1920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 357,
                 
                 P
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b110111; // Expected: {'P': 1430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 358,
                 
                 P
                 , 
                 
                 1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b111111; // Expected: {'P': 2457}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 359,
                 
                 P
                 , 
                 
                 2457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b011110; // Expected: {'P': 1380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 360,
                 
                 P
                 , 
                 
                 1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b010011; // Expected: {'P': 570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 361,
                 
                 P
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b000111; // Expected: {'P': 322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 362,
                 
                 P
                 , 
                 
                 322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b101110; // Expected: {'P': 2024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 363,
                 
                 P
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100000; // Expected: {'P': 608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 364,
                 
                 P
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b110101; // Expected: {'P': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 365,
                 
                 P
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 366,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b110110; // Expected: {'P': 3294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 367,
                 
                 P
                 , 
                 
                 3294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b111110; // Expected: {'P': 434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 368,
                 
                 P
                 , 
                 
                 434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 369,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b111010; // Expected: {'P': 1392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 370,
                 
                 P
                 , 
                 
                 1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b111100; // Expected: {'P': 3660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 371,
                 
                 P
                 , 
                 
                 3660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b110110; // Expected: {'P': 2214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 372,
                 
                 P
                 , 
                 
                 2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 373,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 374,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b000011; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 375,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b000001; // Expected: {'P': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 376,
                 
                 P
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b010110; // Expected: {'P': 484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 377,
                 
                 P
                 , 
                 
                 484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b001001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 378,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000111; // Expected: {'P': 294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 379,
                 
                 P
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b111100; // Expected: {'P': 780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 380,
                 
                 P
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000111; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 381,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b000110; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 382,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b010100; // Expected: {'P': 520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 383,
                 
                 P
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b110111; // Expected: {'P': 2255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 384,
                 
                 P
                 , 
                 
                 2255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b010000; // Expected: {'P': 512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 385,
                 
                 P
                 , 
                 
                 512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b100101; // Expected: {'P': 1073}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 386,
                 
                 P
                 , 
                 
                 1073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b100001; // Expected: {'P': 1683}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 387,
                 
                 P
                 , 
                 
                 1683
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b010110; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 388,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b110000; // Expected: {'P': 1104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 389,
                 
                 P
                 , 
                 
                 1104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b010100; // Expected: {'P': 1220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 390,
                 
                 P
                 , 
                 
                 1220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b111101; // Expected: {'P': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 391,
                 
                 P
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101111; // Expected: {'P': 329}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 392,
                 
                 P
                 , 
                 
                 329
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101101; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 393,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b011100; // Expected: {'P': 812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 394,
                 
                 P
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b010111; // Expected: {'P': 759}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 395,
                 
                 P
                 , 
                 
                 759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b011101; // Expected: {'P': 841}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 396,
                 
                 P
                 , 
                 
                 841
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b110100; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 397,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b011001; // Expected: {'P': 375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 398,
                 
                 P
                 , 
                 
                 375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100111; // Expected: {'P': 351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 399,
                 
                 P
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101011; // Expected: {'P': 1677}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 400,
                 
                 P
                 , 
                 
                 1677
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110001; // Expected: {'P': 2793}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 401,
                 
                 P
                 , 
                 
                 2793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b011000; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 402,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b001101; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 403,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b011101; // Expected: {'P': 1566}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 404,
                 
                 P
                 , 
                 
                 1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b110001; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 405,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 406,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000010; // Expected: {'P': 6}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 407,
                 
                 P
                 , 
                 
                 6
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b101011; // Expected: {'P': 1978}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 408,
                 
                 P
                 , 
                 
                 1978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b010000; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 409,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b010000; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 410,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b001101; // Expected: {'P': 598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 411,
                 
                 P
                 , 
                 
                 598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101101; // Expected: {'P': 2610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 412,
                 
                 P
                 , 
                 
                 2610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b100001; // Expected: {'P': 759}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 413,
                 
                 P
                 , 
                 
                 759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b000011; // Expected: {'P': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 414,
                 
                 P
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b010010; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 415,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b011011; // Expected: {'P': 729}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 416,
                 
                 P
                 , 
                 
                 729
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b101111; // Expected: {'P': 470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 417,
                 
                 P
                 , 
                 
                 470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111110; // Expected: {'P': 2852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 418,
                 
                 P
                 , 
                 
                 2852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b001001; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 419,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b000111; // Expected: {'P': 147}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 420,
                 
                 P
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b100010; // Expected: {'P': 1224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 421,
                 
                 P
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111100; // Expected: {'P': 2280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 422,
                 
                 P
                 , 
                 
                 2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101111; // Expected: {'P': 2585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 423,
                 
                 P
                 , 
                 
                 2585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b011101; // Expected: {'P': 1102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 424,
                 
                 P
                 , 
                 
                 1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b000001; // Expected: {'P': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 425,
                 
                 P
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b101001; // Expected: {'P': 1886}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 426,
                 
                 P
                 , 
                 
                 1886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b110100; // Expected: {'P': 2496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 427,
                 
                 P
                 , 
                 
                 2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b001101; // Expected: {'P': 676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 428,
                 
                 P
                 , 
                 
                 676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 429,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b010010; // Expected: {'P': 972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 430,
                 
                 P
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110000; // Expected: {'P': 2688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 431,
                 
                 P
                 , 
                 
                 2688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b110001; // Expected: {'P': 637}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 432,
                 
                 P
                 , 
                 
                 637
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b000111; // Expected: {'P': 392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 433,
                 
                 P
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b010100; // Expected: {'P': 1100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 434,
                 
                 P
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100010; // Expected: {'P': 1564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 435,
                 
                 P
                 , 
                 
                 1564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b010101; // Expected: {'P': 693}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 436,
                 
                 P
                 , 
                 
                 693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b010101; // Expected: {'P': 1239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 437,
                 
                 P
                 , 
                 
                 1239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b000111; // Expected: {'P': 133}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 438,
                 
                 P
                 , 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b000010; // Expected: {'P': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 439,
                 
                 P
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b101111; // Expected: {'P': 1598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 440,
                 
                 P
                 , 
                 
                 1598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101011; // Expected: {'P': 473}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 441,
                 
                 P
                 , 
                 
                 473
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b110100; // Expected: {'P': 2600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 442,
                 
                 P
                 , 
                 
                 2600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b000001; // Expected: {'P': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 443,
                 
                 P
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b110111; // Expected: {'P': 935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 444,
                 
                 P
                 , 
                 
                 935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b111010; // Expected: {'P': 3190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 445,
                 
                 P
                 , 
                 
                 3190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b010011; // Expected: {'P': 893}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 446,
                 
                 P
                 , 
                 
                 893
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011100; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 447,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b001001; // Expected: {'P': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 448,
                 
                 P
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111111; // Expected: {'P': 3087}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 449,
                 
                 P
                 , 
                 
                 3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b110001; // Expected: {'P': 833}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 450,
                 
                 P
                 , 
                 
                 833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111000; // Expected: {'P': 896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 451,
                 
                 P
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101111; // Expected: {'P': 1833}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 452,
                 
                 P
                 , 
                 
                 1833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b010011; // Expected: {'P': 95}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 453,
                 
                 P
                 , 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b111010; // Expected: {'P': 1624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 454,
                 
                 P
                 , 
                 
                 1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b101001; // Expected: {'P': 1148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 455,
                 
                 P
                 , 
                 
                 1148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b111010; // Expected: {'P': 1856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 456,
                 
                 P
                 , 
                 
                 1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b011001; // Expected: {'P': 1075}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 457,
                 
                 P
                 , 
                 
                 1075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b111010; // Expected: {'P': 1566}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 458,
                 
                 P
                 , 
                 
                 1566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b000101; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 459,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101101; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 460,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b110000; // Expected: {'P': 864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 461,
                 
                 P
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b001000; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 462,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b100001; // Expected: {'P': 1452}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 463,
                 
                 P
                 , 
                 
                 1452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b011000; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 464,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b110111; // Expected: {'P': 1100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 465,
                 
                 P
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111011; // Expected: {'P': 3717}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 466,
                 
                 P
                 , 
                 
                 3717
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b101000; // Expected: {'P': 2280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 467,
                 
                 P
                 , 
                 
                 2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b001011; // Expected: {'P': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 468,
                 
                 P
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b110000; // Expected: {'P': 2640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 469,
                 
                 P
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b010111; // Expected: {'P': 437}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 470,
                 
                 P
                 , 
                 
                 437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100100; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 471,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b010100; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 472,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100100; // Expected: {'P': 684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 473,
                 
                 P
                 , 
                 
                 684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101011; // Expected: {'P': 2709}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 474,
                 
                 P
                 , 
                 
                 2709
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000101; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 475,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b110110; // Expected: {'P': 3348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 476,
                 
                 P
                 , 
                 
                 3348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b100100; // Expected: {'P': 1116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 477,
                 
                 P
                 , 
                 
                 1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010000; // Expected: {'P': 896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 478,
                 
                 P
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100010; // Expected: {'P': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 479,
                 
                 P
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b000010; // Expected: {'P': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 480,
                 
                 P
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b001011; // Expected: {'P': 638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 481,
                 
                 P
                 , 
                 
                 638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010011; // Expected: {'P': 836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 482,
                 
                 P
                 , 
                 
                 836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111001; // Expected: {'P': 912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 483,
                 
                 P
                 , 
                 
                 912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110011; // Expected: {'P': 2703}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 484,
                 
                 P
                 , 
                 
                 2703
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b010001; // Expected: {'P': 782}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 485,
                 
                 P
                 , 
                 
                 782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b010110; // Expected: {'P': 946}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 486,
                 
                 P
                 , 
                 
                 946
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b110001; // Expected: {'P': 2303}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 487,
                 
                 P
                 , 
                 
                 2303
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b100110; // Expected: {'P': 1976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 488,
                 
                 P
                 , 
                 
                 1976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b011100; // Expected: {'P': 980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 489,
                 
                 P
                 , 
                 
                 980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b001111; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 490,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b000100; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 491,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b100101; // Expected: {'P': 74}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 492,
                 
                 P
                 , 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010110; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 493,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b101011; // Expected: {'P': 602}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 494,
                 
                 P
                 , 
                 
                 602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b100110; // Expected: {'P': 2090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 495,
                 
                 P
                 , 
                 
                 2090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b000001; // Expected: {'P': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 496,
                 
                 P
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110100; // Expected: {'P': 2964}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 497,
                 
                 P
                 , 
                 
                 2964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b000101; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 498,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b000110; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 499,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b000111; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 500,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b010100; // Expected: {'P': 780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 501,
                 
                 P
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b100100; // Expected: {'P': 648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 502,
                 
                 P
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111111; // Expected: {'P': 2898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 503,
                 
                 P
                 , 
                 
                 2898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b110001; // Expected: {'P': 2352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 504,
                 
                 P
                 , 
                 
                 2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b001000; // Expected: {'P': 304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 505,
                 
                 P
                 , 
                 
                 304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b100000; // Expected: {'P': 1088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 506,
                 
                 P
                 , 
                 
                 1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b111011; // Expected: {'P': 3422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 507,
                 
                 P
                 , 
                 
                 3422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101000; // Expected: {'P': 2000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 508,
                 
                 P
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b110010; // Expected: {'P': 1350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 509,
                 
                 P
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000010; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 510,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b010001; // Expected: {'P': 867}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 511,
                 
                 P
                 , 
                 
                 867
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b011101; // Expected: {'P': 986}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 512,
                 
                 P
                 , 
                 
                 986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b110001; // Expected: {'P': 1078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 513,
                 
                 P
                 , 
                 
                 1078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011010; // Expected: {'P': 416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 514,
                 
                 P
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b110010; // Expected: {'P': 3050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 515,
                 
                 P
                 , 
                 
                 3050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b011111; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 516,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b101001; // Expected: {'P': 2460}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 517,
                 
                 P
                 , 
                 
                 2460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b100101; // Expected: {'P': 2109}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 518,
                 
                 P
                 , 
                 
                 2109
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b111010; // Expected: {'P': 2610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 519,
                 
                 P
                 , 
                 
                 2610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101101; // Expected: {'P': 2250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 520,
                 
                 P
                 , 
                 
                 2250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b100011; // Expected: {'P': 1400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 521,
                 
                 P
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b101100; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 522,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b001011; // Expected: {'P': 495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 523,
                 
                 P
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b011110; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 524,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b101001; // Expected: {'P': 697}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 525,
                 
                 P
                 , 
                 
                 697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b101110; // Expected: {'P': 368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 526,
                 
                 P
                 , 
                 
                 368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101001; // Expected: {'P': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 527,
                 
                 P
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b010110; // Expected: {'P': 242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 528,
                 
                 P
                 , 
                 
                 242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b110011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 529,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b001001; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 530,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b011011; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 531,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111000; // Expected: {'P': 3528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 532,
                 
                 P
                 , 
                 
                 3528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b111001; // Expected: {'P': 1368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 533,
                 
                 P
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000100; // Expected: {'P': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 534,
                 
                 P
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b101101; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 535,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b001100; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 536,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b001010; // Expected: {'P': 320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 537,
                 
                 P
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b100110; // Expected: {'P': 266}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 538,
                 
                 P
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b001010; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 539,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110100; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 540,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001101; // Expected: {'P': 351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 541,
                 
                 P
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101100; // Expected: {'P': 704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 542,
                 
                 P
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b101100; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 543,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b111111; // Expected: {'P': 3843}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 544,
                 
                 P
                 , 
                 
                 3843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b110111; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 545,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110000; // Expected: {'P': 1488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 546,
                 
                 P
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b000101; // Expected: {'P': 125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 547,
                 
                 P
                 , 
                 
                 125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b111101; // Expected: {'P': 305}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 548,
                 
                 P
                 , 
                 
                 305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 549,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011010; // Expected: {'P': 494}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 550,
                 
                 P
                 , 
                 
                 494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b000100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 551,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b110111; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 552,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101010; // Expected: {'P': 1638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 553,
                 
                 P
                 , 
                 
                 1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 554,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b100110; // Expected: {'P': 950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 555,
                 
                 P
                 , 
                 
                 950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b100101; // Expected: {'P': 1813}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 556,
                 
                 P
                 , 
                 
                 1813
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b000010; // Expected: {'P': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 557,
                 
                 P
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b011101; // Expected: {'P': 638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 558,
                 
                 P
                 , 
                 
                 638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b111101; // Expected: {'P': 1891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 559,
                 
                 P
                 , 
                 
                 1891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110011; // Expected: {'P': 2754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 560,
                 
                 P
                 , 
                 
                 2754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b110101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 561,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b001100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 562,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b010101; // Expected: {'P': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 563,
                 
                 P
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b000011; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 564,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b001001; // Expected: {'P': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 565,
                 
                 P
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b010111; // Expected: {'P': 207}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 566,
                 
                 P
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b100001; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 567,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b000011; // Expected: {'P': 129}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 568,
                 
                 P
                 , 
                 
                 129
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b001000; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 569,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b110101; // Expected: {'P': 371}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 570,
                 
                 P
                 , 
                 
                 371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000101; // Expected: {'P': 295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 571,
                 
                 P
                 , 
                 
                 295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b000110; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 572,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b000111; // Expected: {'P': 175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 573,
                 
                 P
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100010; // Expected: {'P': 476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 574,
                 
                 P
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b010101; // Expected: {'P': 945}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 575,
                 
                 P
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b011011; // Expected: {'P': 567}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 576,
                 
                 P
                 , 
                 
                 567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101111; // Expected: {'P': 517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 577,
                 
                 P
                 , 
                 
                 517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b111101; // Expected: {'P': 854}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 578,
                 
                 P
                 , 
                 
                 854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b011001; // Expected: {'P': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 579,
                 
                 P
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110111; // Expected: {'P': 495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 580,
                 
                 P
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011110; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 581,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b001101; // Expected: {'P': 455}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 582,
                 
                 P
                 , 
                 
                 455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b000100; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 583,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b010110; // Expected: {'P': 704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 584,
                 
                 P
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b111001; // Expected: {'P': 1881}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 585,
                 
                 P
                 , 
                 
                 1881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b101011; // Expected: {'P': 1032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 586,
                 
                 P
                 , 
                 
                 1032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b001000; // Expected: {'P': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 587,
                 
                 P
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b111010; // Expected: {'P': 3306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 588,
                 
                 P
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b111011; // Expected: {'P': 177}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 589,
                 
                 P
                 , 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b111001; // Expected: {'P': 2337}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 590,
                 
                 P
                 , 
                 
                 2337
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b000001; // Expected: {'P': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 591,
                 
                 P
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011001; // Expected: {'P': 1275}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 592,
                 
                 P
                 , 
                 
                 1275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101010; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 593,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b110100; // Expected: {'P': 2184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 594,
                 
                 P
                 , 
                 
                 2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100001; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 595,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110011; // Expected: {'P': 1581}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 596,
                 
                 P
                 , 
                 
                 1581
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000110; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 597,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b011110; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 598,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b101001; // Expected: {'P': 1476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 599,
                 
                 P
                 , 
                 
                 1476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b001111; // Expected: {'P': 675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 600,
                 
                 P
                 , 
                 
                 675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b010101; // Expected: {'P': 1155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 601,
                 
                 P
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 602,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b110000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 603,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b110001; // Expected: {'P': 1862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 604,
                 
                 P
                 , 
                 
                 1862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b000010; // Expected: {'P': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 605,
                 
                 P
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100001; // Expected: {'P': 297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 606,
                 
                 P
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100001; // Expected: {'P': 1485}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 607,
                 
                 P
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101000; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 608,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b001011; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 609,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b100110; // Expected: {'P': 2204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 610,
                 
                 P
                 , 
                 
                 2204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 611,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b110101; // Expected: {'P': 3127}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 612,
                 
                 P
                 , 
                 
                 3127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 613,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b001010; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 614,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b100011; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 615,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b011011; // Expected: {'P': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 616,
                 
                 P
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b011011; // Expected: {'P': 1431}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 617,
                 
                 P
                 , 
                 
                 1431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b111011; // Expected: {'P': 2537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 618,
                 
                 P
                 , 
                 
                 2537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b110000; // Expected: {'P': 768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 619,
                 
                 P
                 , 
                 
                 768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b101000; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 620,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b110100; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 621,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b001111; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 622,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b000100; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 623,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b111010; // Expected: {'P': 2958}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 624,
                 
                 P
                 , 
                 
                 2958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100000; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 625,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b101100; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 626,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b101100; // Expected: {'P': 1584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 627,
                 
                 P
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b011101; // Expected: {'P': 1247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 628,
                 
                 P
                 , 
                 
                 1247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b011001; // Expected: {'P': 1475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 629,
                 
                 P
                 , 
                 
                 1475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b110101; // Expected: {'P': 1431}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 630,
                 
                 P
                 , 
                 
                 1431
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b000001; // Expected: {'P': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 631,
                 
                 P
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b000010; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 632,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b010100; // Expected: {'P': 760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 633,
                 
                 P
                 , 
                 
                 760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b010101; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 634,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b001100; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 635,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b011110; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 636,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b010000; // Expected: {'P': 992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 637,
                 
                 P
                 , 
                 
                 992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101001; // Expected: {'P': 2009}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 638,
                 
                 P
                 , 
                 
                 2009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b111111; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 639,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b001101; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 640,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b111110; // Expected: {'P': 1798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 641,
                 
                 P
                 , 
                 
                 1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110101; // Expected: {'P': 1590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 642,
                 
                 P
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b001000; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 643,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b101100; // Expected: {'P': 2508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 644,
                 
                 P
                 , 
                 
                 2508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b011010; // Expected: {'P': 1352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 645,
                 
                 P
                 , 
                 
                 1352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b100110; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 646,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b011110; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 647,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b101110; // Expected: {'P': 1472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 648,
                 
                 P
                 , 
                 
                 1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b010010; // Expected: {'P': 846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 649,
                 
                 P
                 , 
                 
                 846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 650,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b111001; // Expected: {'P': 1083}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 651,
                 
                 P
                 , 
                 
                 1083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b010100; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 652,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b110010; // Expected: {'P': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 653,
                 
                 P
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b011010; // Expected: {'P': 806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 654,
                 
                 P
                 , 
                 
                 806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b001101; // Expected: {'P': 429}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 655,
                 
                 P
                 , 
                 
                 429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001010; // Expected: {'P': 430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 656,
                 
                 P
                 , 
                 
                 430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b010010; // Expected: {'P': 648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 657,
                 
                 P
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b011001; // Expected: {'P': 575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 658,
                 
                 P
                 , 
                 
                 575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b100000; // Expected: {'P': 640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 659,
                 
                 P
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010110; // Expected: {'P': 1232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 660,
                 
                 P
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b011101; // Expected: {'P': 435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 661,
                 
                 P
                 , 
                 
                 435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001001; // Expected: {'P': 99}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 662,
                 
                 P
                 , 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b001011; // Expected: {'P': 517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 663,
                 
                 P
                 , 
                 
                 517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b110000; // Expected: {'P': 1584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 664,
                 
                 P
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b100001; // Expected: {'P': 2079}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 665,
                 
                 P
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b011010; // Expected: {'P': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 666,
                 
                 P
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b011010; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 667,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011001; // Expected: {'P': 1050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 668,
                 
                 P
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b111001; // Expected: {'P': 2508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 669,
                 
                 P
                 , 
                 
                 2508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b111111; // Expected: {'P': 3717}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 670,
                 
                 P
                 , 
                 
                 3717
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b001011; // Expected: {'P': 572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 671,
                 
                 P
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b110100; // Expected: {'P': 2288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 672,
                 
                 P
                 , 
                 
                 2288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b001100; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 673,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011110; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 674,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101100; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 675,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b110111; // Expected: {'P': 275}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 676,
                 
                 P
                 , 
                 
                 275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b011111; // Expected: {'P': 806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 677,
                 
                 P
                 , 
                 
                 806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b100001; // Expected: {'P': 1914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 678,
                 
                 P
                 , 
                 
                 1914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b011111; // Expected: {'P': 682}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 679,
                 
                 P
                 , 
                 
                 682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100111; // Expected: {'P': 1443}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 680,
                 
                 P
                 , 
                 
                 1443
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b110101; // Expected: {'P': 2650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 681,
                 
                 P
                 , 
                 
                 2650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 682,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010010; // Expected: {'P': 792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 683,
                 
                 P
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b100010; // Expected: {'P': 340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 684,
                 
                 P
                 , 
                 
                 340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b100110; // Expected: {'P': 418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 685,
                 
                 P
                 , 
                 
                 418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100101; // Expected: {'P': 555}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 686,
                 
                 P
                 , 
                 
                 555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b110100; // Expected: {'P': 3068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 687,
                 
                 P
                 , 
                 
                 3068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b110100; // Expected: {'P': 2704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 688,
                 
                 P
                 , 
                 
                 2704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b000010; // Expected: {'P': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 689,
                 
                 P
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101001; // Expected: {'P': 2132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 690,
                 
                 P
                 , 
                 
                 2132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011110; // Expected: {'P': 1410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 691,
                 
                 P
                 , 
                 
                 1410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b111000; // Expected: {'P': 2800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 692,
                 
                 P
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b001011; // Expected: {'P': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 693,
                 
                 P
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b100010; // Expected: {'P': 1870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 694,
                 
                 P
                 , 
                 
                 1870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b000001; // Expected: {'P': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 695,
                 
                 P
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b111011; // Expected: {'P': 1770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 696,
                 
                 P
                 , 
                 
                 1770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b010001; // Expected: {'P': 459}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 697,
                 
                 P
                 , 
                 
                 459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b010011; // Expected: {'P': 266}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 698,
                 
                 P
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b000011; // Expected: {'P': 153}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 699,
                 
                 P
                 , 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b010100; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 700,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b010001; // Expected: {'P': 544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 701,
                 
                 P
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b011001; // Expected: {'P': 875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 702,
                 
                 P
                 , 
                 
                 875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000110; // Expected: {'P': 354}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 703,
                 
                 P
                 , 
                 
                 354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b101001; // Expected: {'P': 1394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 704,
                 
                 P
                 , 
                 
                 1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b110000; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 705,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110010; // Expected: {'P': 2800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 706,
                 
                 P
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b111000; // Expected: {'P': 1624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 707,
                 
                 P
                 , 
                 
                 1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b100011; // Expected: {'P': 875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 708,
                 
                 P
                 , 
                 
                 875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101001; // Expected: {'P': 451}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 709,
                 
                 P
                 , 
                 
                 451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101101; // Expected: {'P': 495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 710,
                 
                 P
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b000101; // Expected: {'P': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 711,
                 
                 P
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b110001; // Expected: {'P': 2156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 712,
                 
                 P
                 , 
                 
                 2156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b100100; // Expected: {'P': 1944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 713,
                 
                 P
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b111000; // Expected: {'P': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 714,
                 
                 P
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b110001; // Expected: {'P': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 715,
                 
                 P
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b101111; // Expected: {'P': 1222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 716,
                 
                 P
                 , 
                 
                 1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b000111; // Expected: {'P': 259}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 717,
                 
                 P
                 , 
                 
                 259
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b001111; // Expected: {'P': 105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 718,
                 
                 P
                 , 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b101100; // Expected: {'P': 1012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 719,
                 
                 P
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b111000; // Expected: {'P': 2184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 720,
                 
                 P
                 , 
                 
                 2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001000; // Expected: {'P': 344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 721,
                 
                 P
                 , 
                 
                 344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b011100; // Expected: {'P': 784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 722,
                 
                 P
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b110001; // Expected: {'P': 3087}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 723,
                 
                 P
                 , 
                 
                 3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b011010; // Expected: {'P': 1196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 724,
                 
                 P
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b101101; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 725,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b100000; // Expected: {'P': 1952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 726,
                 
                 P
                 , 
                 
                 1952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b010100; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 727,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b100111; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 728,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b111010; // Expected: {'P': 2726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 729,
                 
                 P
                 , 
                 
                 2726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010111; // Expected: {'P': 1012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 730,
                 
                 P
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111111; // Expected: {'P': 567}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 731,
                 
                 P
                 , 
                 
                 567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b111100; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 732,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b111011; // Expected: {'P': 1357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 733,
                 
                 P
                 , 
                 
                 1357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b001001; // Expected: {'P': 441}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 734,
                 
                 P
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b110001; // Expected: {'P': 294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 735,
                 
                 P
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b110111; // Expected: {'P': 1375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 736,
                 
                 P
                 , 
                 
                 1375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010110; // Expected: {'P': 968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 737,
                 
                 P
                 , 
                 
                 968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b011101; // Expected: {'P': 203}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 738,
                 
                 P
                 , 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b000111; // Expected: {'P': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 739,
                 
                 P
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011100; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 740,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b000011; // Expected: {'P': 123}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 741,
                 
                 P
                 , 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b011111; // Expected: {'P': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 742,
                 
                 P
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b100001; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 743,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b011111; // Expected: {'P': 403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 744,
                 
                 P
                 , 
                 
                 403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b110001; // Expected: {'P': 1323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 745,
                 
                 P
                 , 
                 
                 1323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b101010; // Expected: {'P': 2352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 746,
                 
                 P
                 , 
                 
                 2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010101; // Expected: {'P': 651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 747,
                 
                 P
                 , 
                 
                 651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b001101; // Expected: {'P': 754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 748,
                 
                 P
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100101; // Expected: {'P': 518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 749,
                 
                 P
                 , 
                 
                 518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111000; // Expected: {'P': 2128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 750,
                 
                 P
                 , 
                 
                 2128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b110111; // Expected: {'P': 2585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 751,
                 
                 P
                 , 
                 
                 2585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101101; // Expected: {'P': 2295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 752,
                 
                 P
                 , 
                 
                 2295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b001101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 753,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101000; // Expected: {'P': 1960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 754,
                 
                 P
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b001001; // Expected: {'P': 423}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 755,
                 
                 P
                 , 
                 
                 423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b001100; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 756,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b101001; // Expected: {'P': 861}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 757,
                 
                 P
                 , 
                 
                 861
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b101111; // Expected: {'P': 1880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 758,
                 
                 P
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b111000; // Expected: {'P': 448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 759,
                 
                 P
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111000; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 760,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b101001; // Expected: {'P': 2337}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 761,
                 
                 P
                 , 
                 
                 2337
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000011; // Expected: {'P': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 762,
                 
                 P
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110101; // Expected: {'P': 159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 763,
                 
                 P
                 , 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b000110; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 764,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b010111; // Expected: {'P': 460}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 765,
                 
                 P
                 , 
                 
                 460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b000111; // Expected: {'P': 287}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 766,
                 
                 P
                 , 
                 
                 287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b101011; // Expected: {'P': 344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 767,
                 
                 P
                 , 
                 
                 344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b010101; // Expected: {'P': 1071}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 768,
                 
                 P
                 , 
                 
                 1071
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b111101; // Expected: {'P': 3355}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 769,
                 
                 P
                 , 
                 
                 3355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b010100; // Expected: {'P': 320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 770,
                 
                 P
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b111100; // Expected: {'P': 1140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 771,
                 
                 P
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b110100; // Expected: {'P': 988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 772,
                 
                 P
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b100011; // Expected: {'P': 245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 773,
                 
                 P
                 , 
                 
                 245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b010111; // Expected: {'P': 552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 774,
                 
                 P
                 , 
                 
                 552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b101000; // Expected: {'P': 1280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 775,
                 
                 P
                 , 
                 
                 1280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b101001; // Expected: {'P': 123}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 776,
                 
                 P
                 , 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b100101; // Expected: {'P': 111}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 777,
                 
                 P
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110110; // Expected: {'P': 3078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 778,
                 
                 P
                 , 
                 
                 3078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b111011; // Expected: {'P': 1475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 779,
                 
                 P
                 , 
                 
                 1475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b001010; // Expected: {'P': 490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 780,
                 
                 P
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101100; // Expected: {'P': 2244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 781,
                 
                 P
                 , 
                 
                 2244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b001011; // Expected: {'P': 561}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 782,
                 
                 P
                 , 
                 
                 561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b011111; // Expected: {'P': 651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 783,
                 
                 P
                 , 
                 
                 651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b010110; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 784,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010001; // Expected: {'P': 102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 785,
                 
                 P
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101010; // Expected: {'P': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 786,
                 
                 P
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b110110; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 787,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b110001; // Expected: {'P': 588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 788,
                 
                 P
                 , 
                 
                 588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b000100; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 789,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b101011; // Expected: {'P': 387}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 790,
                 
                 P
                 , 
                 
                 387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b001001; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 791,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b001001; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 792,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010010; // Expected: {'P': 738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 793,
                 
                 P
                 , 
                 
                 738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b101101; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 794,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b100010; // Expected: {'P': 1734}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 795,
                 
                 P
                 , 
                 
                 1734
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b101011; // Expected: {'P': 903}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 796,
                 
                 P
                 , 
                 
                 903
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011110; // Expected: {'P': 570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 797,
                 
                 P
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b001111; // Expected: {'P': 765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 798,
                 
                 P
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b001000; // Expected: {'P': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 799,
                 
                 P
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b111001; // Expected: {'P': 741}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 800,
                 
                 P
                 , 
                 
                 741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b011101; // Expected: {'P': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 801,
                 
                 P
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b011101; // Expected: {'P': 1798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 802,
                 
                 P
                 , 
                 
                 1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111001; // Expected: {'P': 513}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 803,
                 
                 P
                 , 
                 
                 513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001000; // Expected: {'P': 488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 804,
                 
                 P
                 , 
                 
                 488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b100000; // Expected: {'P': 512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 805,
                 
                 P
                 , 
                 
                 512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b110101; // Expected: {'P': 1007}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 806,
                 
                 P
                 , 
                 
                 1007
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b000001; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 807,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b001110; // Expected: {'P': 574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 808,
                 
                 P
                 , 
                 
                 574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b010101; // Expected: {'P': 546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 809,
                 
                 P
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b101110; // Expected: {'P': 1242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 810,
                 
                 P
                 , 
                 
                 1242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b011101; // Expected: {'P': 1044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 811,
                 
                 P
                 , 
                 
                 1044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b011001; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 812,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b100011; // Expected: {'P': 1645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 813,
                 
                 P
                 , 
                 
                 1645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b000011; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 814,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110110; // Expected: {'P': 3024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 815,
                 
                 P
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101011; // Expected: {'P': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 816,
                 
                 P
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b000011; // Expected: {'P': 111}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 817,
                 
                 P
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b111111; // Expected: {'P': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 818,
                 
                 P
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b100000; // Expected: {'P': 1984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 819,
                 
                 P
                 , 
                 
                 1984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b111011; // Expected: {'P': 2596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 820,
                 
                 P
                 , 
                 
                 2596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010101; // Expected: {'P': 273}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 821,
                 
                 P
                 , 
                 
                 273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b000111; // Expected: {'P': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 822,
                 
                 P
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b011101; // Expected: {'P': 812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 823,
                 
                 P
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b110011; // Expected: {'P': 1938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 824,
                 
                 P
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b100100; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 825,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b101001; // Expected: {'P': 533}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 826,
                 
                 P
                 , 
                 
                 533
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b011110; // Expected: {'P': 1590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 827,
                 
                 P
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b111001; // Expected: {'P': 1482}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 828,
                 
                 P
                 , 
                 
                 1482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b110101; // Expected: {'P': 689}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 829,
                 
                 P
                 , 
                 
                 689
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b101010; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 830,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b000100; // Expected: {'P': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 831,
                 
                 P
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b110110; // Expected: {'P': 702}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 832,
                 
                 P
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110101; // Expected: {'P': 2862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 833,
                 
                 P
                 , 
                 
                 2862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b111100; // Expected: {'P': 3360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 834,
                 
                 P
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b100000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 835,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b001011; // Expected: {'P': 363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 836,
                 
                 P
                 , 
                 
                 363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b011011; // Expected: {'P': 1620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 837,
                 
                 P
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b011011; // Expected: {'P': 1593}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 838,
                 
                 P
                 , 
                 
                 1593
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100101; // Expected: {'P': 333}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 839,
                 
                 P
                 , 
                 
                 333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 840,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b100110; // Expected: {'P': 2318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 841,
                 
                 P
                 , 
                 
                 2318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b001110; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 842,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b001010; // Expected: {'P': 510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 843,
                 
                 P
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100111; // Expected: {'P': 1638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 844,
                 
                 P
                 , 
                 
                 1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b111101; // Expected: {'P': 671}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 845,
                 
                 P
                 , 
                 
                 671
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b010011; // Expected: {'P': 399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 846,
                 
                 P
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000010; // Expected: {'P': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 847,
                 
                 P
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011111; // Expected: {'P': 1953}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 848,
                 
                 P
                 , 
                 
                 1953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b011101; // Expected: {'P': 1769}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 849,
                 
                 P
                 , 
                 
                 1769
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b001001; // Expected: {'P': 486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 850,
                 
                 P
                 , 
                 
                 486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b111000; // Expected: {'P': 2912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 851,
                 
                 P
                 , 
                 
                 2912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b001010; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 852,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b111100; // Expected: {'P': 3540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 853,
                 
                 P
                 , 
                 
                 3540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b110100; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 854,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b001101; // Expected: {'P': 689}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 855,
                 
                 P
                 , 
                 
                 689
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b101110; // Expected: {'P': 2438}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 856,
                 
                 P
                 , 
                 
                 2438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101011; // Expected: {'P': 301}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 857,
                 
                 P
                 , 
                 
                 301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b010010; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 858,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b100100; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 859,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101110; // Expected: {'P': 736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 860,
                 
                 P
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b101000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 861,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101010; // Expected: {'P': 2436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 862,
                 
                 P
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b000101; // Expected: {'P': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 863,
                 
                 P
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b010100; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 864,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b100101; // Expected: {'P': 592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 865,
                 
                 P
                 , 
                 
                 592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001100; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 866,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b110111; // Expected: {'P': 2365}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 867,
                 
                 P
                 , 
                 
                 2365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 868,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000001; // Expected: {'P': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 869,
                 
                 P
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b010011; // Expected: {'P': 361}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 870,
                 
                 P
                 , 
                 
                 361
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b011001; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 871,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b100100; // Expected: {'P': 1548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 872,
                 
                 P
                 , 
                 
                 1548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101001; // Expected: {'P': 287}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 873,
                 
                 P
                 , 
                 
                 287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b001010; // Expected: {'P': 410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 874,
                 
                 P
                 , 
                 
                 410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b000111; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 875,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b001111; // Expected: {'P': 570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 876,
                 
                 P
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b000100; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 877,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000101; // Expected: {'P': 175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 878,
                 
                 P
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b111001; // Expected: {'P': 627}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 879,
                 
                 P
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b001000; // Expected: {'P': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 880,
                 
                 P
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b111111; // Expected: {'P': 1764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 881,
                 
                 P
                 , 
                 
                 1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001101; // Expected: {'P': 559}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 882,
                 
                 P
                 , 
                 
                 559
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b010010; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 883,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110001; // Expected: {'P': 490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 884,
                 
                 P
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100110; // Expected: {'P': 532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 885,
                 
                 P
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b000110; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 886,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b110111; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 887,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b000001; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 888,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b000001; // Expected: {'P': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 889,
                 
                 P
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b001010; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 890,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 891,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 892,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b010110; // Expected: {'P': 1012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 893,
                 
                 P
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b001100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 894,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b101001; // Expected: {'P': 574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 895,
                 
                 P
                 , 
                 
                 574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b011001; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 896,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b000110; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 897,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b111111; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 898,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b110101; // Expected: {'P': 1060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 899,
                 
                 P
                 , 
                 
                 1060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110000; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 900,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b110111; // Expected: {'P': 2420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 901,
                 
                 P
                 , 
                 
                 2420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b101100; // Expected: {'P': 352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 902,
                 
                 P
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b110101; // Expected: {'P': 1325}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 903,
                 
                 P
                 , 
                 
                 1325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000101; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 904,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b110110; // Expected: {'P': 810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 905,
                 
                 P
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b001110; // Expected: {'P': 728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 906,
                 
                 P
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b001111; // Expected: {'P': 690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 907,
                 
                 P
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100010; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 908,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b010100; // Expected: {'P': 340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 909,
                 
                 P
                 , 
                 
                 340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b100000; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 910,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b011111; // Expected: {'P': 1798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 911,
                 
                 P
                 , 
                 
                 1798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b010110; // Expected: {'P': 1078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 912,
                 
                 P
                 , 
                 
                 1078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000110; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 913,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b011110; // Expected: {'P': 510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 914,
                 
                 P
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b101000; // Expected: {'P': 1720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 915,
                 
                 P
                 , 
                 
                 1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000101; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 916,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100011; // Expected: {'P': 1435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 917,
                 
                 P
                 , 
                 
                 1435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b100010; // Expected: {'P': 680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 918,
                 
                 P
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b110110; // Expected: {'P': 1998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 919,
                 
                 P
                 , 
                 
                 1998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b110110; // Expected: {'P': 648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 920,
                 
                 P
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101100; // Expected: {'P': 2552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 921,
                 
                 P
                 , 
                 
                 2552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b001101; // Expected: {'P': 715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 922,
                 
                 P
                 , 
                 
                 715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b010101; // Expected: {'P': 1302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 923,
                 
                 P
                 , 
                 
                 1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b101011; // Expected: {'P': 86}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 924,
                 
                 P
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b100010; // Expected: {'P': 1632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 925,
                 
                 P
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b101000; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 926,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b010100; // Expected: {'P': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 927,
                 
                 P
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b111001; // Expected: {'P': 1539}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 928,
                 
                 P
                 , 
                 
                 1539
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b111101; // Expected: {'P': 1403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 929,
                 
                 P
                 , 
                 
                 1403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b101111; // Expected: {'P': 564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 930,
                 
                 P
                 , 
                 
                 564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b001001; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 931,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110001; // Expected: {'P': 2597}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 932,
                 
                 P
                 , 
                 
                 2597
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b000001; // Expected: {'P': 13}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 933,
                 
                 P
                 , 
                 
                 13
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101101; // Expected: {'P': 2475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 934,
                 
                 P
                 , 
                 
                 2475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b000111; // Expected: {'P': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 935,
                 
                 P
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b001001; // Expected: {'P': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 936,
                 
                 P
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b101110; // Expected: {'P': 2116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 937,
                 
                 P
                 , 
                 
                 2116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101010; // Expected: {'P': 2184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 938,
                 
                 P
                 , 
                 
                 2184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000110; // Expected: {'P': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 939,
                 
                 P
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b111001; // Expected: {'P': 3306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 940,
                 
                 P
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b110010; // Expected: {'P': 2750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 941,
                 
                 P
                 , 
                 
                 2750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b000011; // Expected: {'P': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 942,
                 
                 P
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b101000; // Expected: {'P': 2440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 943,
                 
                 P
                 , 
                 
                 2440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b111111; // Expected: {'P': 2079}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 944,
                 
                 P
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001001; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 945,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b100011; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 946,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b000010; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 947,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110011; // Expected: {'P': 1989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 948,
                 
                 P
                 , 
                 
                 1989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100011; // Expected: {'P': 665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 949,
                 
                 P
                 , 
                 
                 665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b101110; // Expected: {'P': 1932}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 950,
                 
                 P
                 , 
                 
                 1932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b010101; // Expected: {'P': 1197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 951,
                 
                 P
                 , 
                 
                 1197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b111011; // Expected: {'P': 2065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 952,
                 
                 P
                 , 
                 
                 2065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001010; // Expected: {'P': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 953,
                 
                 P
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b111100; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 954,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b100011; // Expected: {'P': 2030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 955,
                 
                 P
                 , 
                 
                 2030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b110111; // Expected: {'P': 2695}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 956,
                 
                 P
                 , 
                 
                 2695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011001; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 957,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b110011; // Expected: {'P': 51}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 958,
                 
                 P
                 , 
                 
                 51
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110110; // Expected: {'P': 2862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 959,
                 
                 P
                 , 
                 
                 2862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b101000; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 960,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000111; // Expected: {'P': 427}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 961,
                 
                 P
                 , 
                 
                 427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b101000; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 962,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000111; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 963,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b101101; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 964,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b001011; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 965,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b101001; // Expected: {'P': 1722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 966,
                 
                 P
                 , 
                 
                 1722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011011; // Expected: {'P': 1269}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 967,
                 
                 P
                 , 
                 
                 1269
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b000001; // Expected: {'P': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 968,
                 
                 P
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b110010; // Expected: {'P': 1750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 969,
                 
                 P
                 , 
                 
                 1750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b011110; // Expected: {'P': 1860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 970,
                 
                 P
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000010; // Expected: {'P': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 971,
                 
                 P
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 972,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b011010; // Expected: {'P': 728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 973,
                 
                 P
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b101010; // Expected: {'P': 588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 974,
                 
                 P
                 , 
                 
                 588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b100011; // Expected: {'P': 1190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 975,
                 
                 P
                 , 
                 
                 1190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b110111; // Expected: {'P': 3300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 976,
                 
                 P
                 , 
                 
                 3300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b111111; // Expected: {'P': 2583}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 977,
                 
                 P
                 , 
                 
                 2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b010110; // Expected: {'P': 572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 978,
                 
                 P
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001011; // Expected: {'P': 550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 979,
                 
                 P
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b000100; // Expected: {'P': 64}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 980,
                 
                 P
                 , 
                 
                 64
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100000; // Expected: {'P': 448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 981,
                 
                 P
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b101011; // Expected: {'P': 1806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 982,
                 
                 P
                 , 
                 
                 1806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b011110; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 983,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b111110; // Expected: {'P': 3472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 984,
                 
                 P
                 , 
                 
                 3472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010101; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 985,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b000010; // Expected: {'P': 86}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 986,
                 
                 P
                 , 
                 
                 86
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b010100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 987,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000010; // Expected: {'P': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 988,
                 
                 P
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b001011; // Expected: {'P': 627}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 989,
                 
                 P
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101010; // Expected: {'P': 294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 990,
                 
                 P
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b111010; // Expected: {'P': 754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 991,
                 
                 P
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b000100; // Expected: {'P': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 992,
                 
                 P
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b011010; // Expected: {'P': 1560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 993,
                 
                 P
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b001110; // Expected: {'P': 784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 994,
                 
                 P
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b001100; // Expected: {'P': 708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 995,
                 
                 P
                 , 
                 
                 708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b011100; // Expected: {'P': 616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 996,
                 
                 P
                 , 
                 
                 616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b011100; // Expected: {'P': 1708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 997,
                 
                 P
                 , 
                 
                 1708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000111; // Expected: {'P': 413}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 998,
                 
                 P
                 , 
                 
                 413
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b001010; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 999,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101100; // Expected: {'P': 2420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1000,
                 
                 P
                 , 
                 
                 2420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b101110; // Expected: {'P': 874}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1001,
                 
                 P
                 , 
                 
                 874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b011110; // Expected: {'P': 1710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1002,
                 
                 P
                 , 
                 
                 1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000010; // Expected: {'P': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1003,
                 
                 P
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b011001; // Expected: {'P': 1350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1004,
                 
                 P
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000110; // Expected: {'P': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1005,
                 
                 P
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000001; // Expected: {'P': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1006,
                 
                 P
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b001111; // Expected: {'P': 885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1007,
                 
                 P
                 , 
                 
                 885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110000; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1008,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b001110; // Expected: {'P': 686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1009,
                 
                 P
                 , 
                 
                 686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001111; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1010,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b010111; // Expected: {'P': 391}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1011,
                 
                 P
                 , 
                 
                 391
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b100001; // Expected: {'P': 1716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1012,
                 
                 P
                 , 
                 
                 1716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b011010; // Expected: {'P': 1508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1013,
                 
                 P
                 , 
                 
                 1508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b010010; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1014,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101000; // Expected: {'P': 1560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1015,
                 
                 P
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b011001; // Expected: {'P': 525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1016,
                 
                 P
                 , 
                 
                 525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b111001; // Expected: {'P': 3135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1017,
                 
                 P
                 , 
                 
                 3135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b011010; // Expected: {'P': 1586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1018,
                 
                 P
                 , 
                 
                 1586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b101001; // Expected: {'P': 1681}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1019,
                 
                 P
                 , 
                 
                 1681
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b001111; // Expected: {'P': 285}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1020,
                 
                 P
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b101100; // Expected: {'P': 748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1021,
                 
                 P
                 , 
                 
                 748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b001110; // Expected: {'P': 406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1022,
                 
                 P
                 , 
                 
                 406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b110100; // Expected: {'P': 1820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1023,
                 
                 P
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b100000; // Expected: {'P': 2016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1024,
                 
                 P
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b010001; // Expected: {'P': 901}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1025,
                 
                 P
                 , 
                 
                 901
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b001101; // Expected: {'P': 65}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1026,
                 
                 P
                 , 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101101; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1027,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100101; // Expected: {'P': 1369}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1028,
                 
                 P
                 , 
                 
                 1369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b100100; // Expected: {'P': 2232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1029,
                 
                 P
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b001010; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1030,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b101111; // Expected: {'P': 1363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1031,
                 
                 P
                 , 
                 
                 1363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b101101; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1032,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b001110; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1033,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b110100; // Expected: {'P': 572}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1034,
                 
                 P
                 , 
                 
                 572
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b011010; // Expected: {'P': 962}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1035,
                 
                 P
                 , 
                 
                 962
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b000111; // Expected: {'P': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1036,
                 
                 P
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b111011; // Expected: {'P': 472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1037,
                 
                 P
                 , 
                 
                 472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b111010; // Expected: {'P': 2378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1038,
                 
                 P
                 , 
                 
                 2378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b001000; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1039,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b111000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1040,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100110; // Expected: {'P': 342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1041,
                 
                 P
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b111100; // Expected: {'P': 3420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1042,
                 
                 P
                 , 
                 
                 3420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b110010; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1043,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001001; // Expected: {'P': 387}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1044,
                 
                 P
                 , 
                 
                 387
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b111111; // Expected: {'P': 1386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1045,
                 
                 P
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b110111; // Expected: {'P': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1046,
                 
                 P
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b001011; // Expected: {'P': 583}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1047,
                 
                 P
                 , 
                 
                 583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1048,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b100000; // Expected: {'P': 1568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1049,
                 
                 P
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b010111; // Expected: {'P': 345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1050,
                 
                 P
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b000011; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1051,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b100101; // Expected: {'P': 1961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1052,
                 
                 P
                 , 
                 
                 1961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b101000; // Expected: {'P': 2400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1053,
                 
                 P
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101111; // Expected: {'P': 2303}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1054,
                 
                 P
                 , 
                 
                 2303
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b100000; // Expected: {'P': 1792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1055,
                 
                 P
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b011010; // Expected: {'P': 1482}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1056,
                 
                 P
                 , 
                 
                 1482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b101010; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1057,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100100; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1058,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b010010; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1059,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b110111; // Expected: {'P': 2090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1060,
                 
                 P
                 , 
                 
                 2090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b100100; // Expected: {'P': 612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1061,
                 
                 P
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b111000; // Expected: {'P': 1400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1062,
                 
                 P
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001011; // Expected: {'P': 297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1063,
                 
                 P
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b101100; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1064,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100001; // Expected: {'P': 1386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1065,
                 
                 P
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b010001; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1066,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100011; // Expected: {'P': 945}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1067,
                 
                 P
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b010101; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1068,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b100011; // Expected: {'P': 1960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1069,
                 
                 P
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b000001; // Expected: {'P': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1070,
                 
                 P
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b010000; // Expected: {'P': 272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1071,
                 
                 P
                 , 
                 
                 272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101011; // Expected: {'P': 2494}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1072,
                 
                 P
                 , 
                 
                 2494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b011010; // Expected: {'P': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1073,
                 
                 P
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100011; // Expected: {'P': 490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1074,
                 
                 P
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b111010; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1075,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b010000; // Expected: {'P': 304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1076,
                 
                 P
                 , 
                 
                 304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b100100; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1077,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b100100; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1078,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b011010; // Expected: {'P': 910}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1079,
                 
                 P
                 , 
                 
                 910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b111011; // Expected: {'P': 3009}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1080,
                 
                 P
                 , 
                 
                 3009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b100010; // Expected: {'P': 1088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1081,
                 
                 P
                 , 
                 
                 1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b010101; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1082,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011101; // Expected: {'P': 1479}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1083,
                 
                 P
                 , 
                 
                 1479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101100; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1084,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b100111; // Expected: {'P': 975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1085,
                 
                 P
                 , 
                 
                 975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b110011; // Expected: {'P': 1071}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1086,
                 
                 P
                 , 
                 
                 1071
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b011001; // Expected: {'P': 650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1087,
                 
                 P
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b100111; // Expected: {'P': 1833}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1088,
                 
                 P
                 , 
                 
                 1833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b011001; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1089,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101101; // Expected: {'P': 1755}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1090,
                 
                 P
                 , 
                 
                 1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001010; // Expected: {'P': 340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1091,
                 
                 P
                 , 
                 
                 340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011010; // Expected: {'P': 1638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1092,
                 
                 P
                 , 
                 
                 1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001111; // Expected: {'P': 645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1093,
                 
                 P
                 , 
                 
                 645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b011011; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1094,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b001110; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1095,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b011111; // Expected: {'P': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1096,
                 
                 P
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b111000; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1097,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b010011; // Expected: {'P': 931}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1098,
                 
                 P
                 , 
                 
                 931
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111000; // Expected: {'P': 3360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1099,
                 
                 P
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b100110; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1100,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110100; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1101,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b111111; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1102,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b111101; // Expected: {'P': 1220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1103,
                 
                 P
                 , 
                 
                 1220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011101; // Expected: {'P': 696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1104,
                 
                 P
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b011001; // Expected: {'P': 825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1105,
                 
                 P
                 , 
                 
                 825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b101000; // Expected: {'P': 1360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1106,
                 
                 P
                 , 
                 
                 1360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b110011; // Expected: {'P': 2397}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1107,
                 
                 P
                 , 
                 
                 2397
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b010000; // Expected: {'P': 864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1108,
                 
                 P
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b110011; // Expected: {'P': 2448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1109,
                 
                 P
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001001; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1110,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b010010; // Expected: {'P': 342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1111,
                 
                 P
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100000; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1112,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101101; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1113,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b110010; // Expected: {'P': 2900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1114,
                 
                 P
                 , 
                 
                 2900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b100001; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1115,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b001011; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1116,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b101110; // Expected: {'P': 2760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1117,
                 
                 P
                 , 
                 
                 2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b110010; // Expected: {'P': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1118,
                 
                 P
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b010111; // Expected: {'P': 69}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1119,
                 
                 P
                 , 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b010110; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1120,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101110; // Expected: {'P': 1610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1121,
                 
                 P
                 , 
                 
                 1610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b100010; // Expected: {'P': 816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1122,
                 
                 P
                 , 
                 
                 816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b010100; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1123,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000011; // Expected: {'P': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1124,
                 
                 P
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b011110; // Expected: {'P': 1560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1125,
                 
                 P
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b010001; // Expected: {'P': 374}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1126,
                 
                 P
                 , 
                 
                 374
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b111100; // Expected: {'P': 2880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1127,
                 
                 P
                 , 
                 
                 2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b011011; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1128,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b001001; // Expected: {'P': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1129,
                 
                 P
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b101010; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1130,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b011101; // Expected: {'P': 377}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1131,
                 
                 P
                 , 
                 
                 377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011010; // Expected: {'P': 1326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1132,
                 
                 P
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100110; // Expected: {'P': 570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1133,
                 
                 P
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b111111; // Expected: {'P': 2772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1134,
                 
                 P
                 , 
                 
                 2772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b001100; // Expected: {'P': 552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1135,
                 
                 P
                 , 
                 
                 552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b001101; // Expected: {'P': 325}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1136,
                 
                 P
                 , 
                 
                 325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b011000; // Expected: {'P': 1296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1137,
                 
                 P
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b110111; // Expected: {'P': 1265}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1138,
                 
                 P
                 , 
                 
                 1265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b010000; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1139,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b011001; // Expected: {'P': 850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1140,
                 
                 P
                 , 
                 
                 850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101011; // Expected: {'P': 2150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1141,
                 
                 P
                 , 
                 
                 2150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010000; // Expected: {'P': 496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1142,
                 
                 P
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b110101; // Expected: {'P': 1749}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1143,
                 
                 P
                 , 
                 
                 1749
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101110; // Expected: {'P': 2668}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1144,
                 
                 P
                 , 
                 
                 2668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b100010; // Expected: {'P': 1326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1145,
                 
                 P
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101101; // Expected: {'P': 2835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1146,
                 
                 P
                 , 
                 
                 2835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b100111; // Expected: {'P': 1911}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1147,
                 
                 P
                 , 
                 
                 1911
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b100111; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1148,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b101101; // Expected: {'P': 2655}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1149,
                 
                 P
                 , 
                 
                 2655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b010011; // Expected: {'P': 380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1150,
                 
                 P
                 , 
                 
                 380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b111101; // Expected: {'P': 1647}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1151,
                 
                 P
                 , 
                 
                 1647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b000110; // Expected: {'P': 258}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1152,
                 
                 P
                 , 
                 
                 258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101011; // Expected: {'P': 2193}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1153,
                 
                 P
                 , 
                 
                 2193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b101111; // Expected: {'P': 846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1154,
                 
                 P
                 , 
                 
                 846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b010000; // Expected: {'P': 800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1155,
                 
                 P
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b111111; // Expected: {'P': 2268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1156,
                 
                 P
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b001000; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1157,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b010100; // Expected: {'P': 920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1158,
                 
                 P
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b011110; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1159,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b110101; // Expected: {'P': 3339}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1160,
                 
                 P
                 , 
                 
                 3339
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b111111; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1161,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b000011; // Expected: {'P': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1162,
                 
                 P
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b100000; // Expected: {'P': 768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1163,
                 
                 P
                 , 
                 
                 768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b010001; // Expected: {'P': 629}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1164,
                 
                 P
                 , 
                 
                 629
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b100000; // Expected: {'P': 704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1165,
                 
                 P
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b111110; // Expected: {'P': 2046}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1166,
                 
                 P
                 , 
                 
                 2046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b010010; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1167,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b001011; // Expected: {'P': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1168,
                 
                 P
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b010010; // Expected: {'P': 954}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1169,
                 
                 P
                 , 
                 
                 954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b011101; // Expected: {'P': 493}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1170,
                 
                 P
                 , 
                 
                 493
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b101011; // Expected: {'P': 1462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1171,
                 
                 P
                 , 
                 
                 1462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b011100; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1172,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b111010; // Expected: {'P': 3364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1173,
                 
                 P
                 , 
                 
                 3364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b000010; // Expected: {'P': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1174,
                 
                 P
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b000011; // Expected: {'P': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1175,
                 
                 P
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b010101; // Expected: {'P': 1218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1176,
                 
                 P
                 , 
                 
                 1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000101; // Expected: {'P': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1177,
                 
                 P
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b101111; // Expected: {'P': 1974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1178,
                 
                 P
                 , 
                 
                 1974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b100100; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1179,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1180,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101000; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1181,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b111101; // Expected: {'P': 427}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1182,
                 
                 P
                 , 
                 
                 427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b001010; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1183,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b110100; // Expected: {'P': 1352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1184,
                 
                 P
                 , 
                 
                 1352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b111001; // Expected: {'P': 2964}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1185,
                 
                 P
                 , 
                 
                 2964
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b001000; // Expected: {'P': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1186,
                 
                 P
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110111; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1187,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b111001; // Expected: {'P': 399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1188,
                 
                 P
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111100; // Expected: {'P': 2940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1189,
                 
                 P
                 , 
                 
                 2940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110100; // Expected: {'P': 520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1190,
                 
                 P
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b100001; // Expected: {'P': 561}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1191,
                 
                 P
                 , 
                 
                 561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b101010; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1192,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001010; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1193,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b111011; // Expected: {'P': 295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1194,
                 
                 P
                 , 
                 
                 295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b111111; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1195,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b001000; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1196,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b100110; // Expected: {'P': 1900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1197,
                 
                 P
                 , 
                 
                 1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b000111; // Expected: {'P': 357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1198,
                 
                 P
                 , 
                 
                 357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b001001; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1199,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001100; // Expected: {'P': 576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1200,
                 
                 P
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b110101; // Expected: {'P': 2226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1201,
                 
                 P
                 , 
                 
                 2226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101000; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1202,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011011; // Expected: {'P': 513}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1203,
                 
                 P
                 , 
                 
                 513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b001001; // Expected: {'P': 117}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1204,
                 
                 P
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b110111; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1205,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b011011; // Expected: {'P': 1242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1206,
                 
                 P
                 , 
                 
                 1242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b111000; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1207,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b101000; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1208,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b111010; // Expected: {'P': 3248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1209,
                 
                 P
                 , 
                 
                 3248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111110; // Expected: {'P': 992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1210,
                 
                 P
                 , 
                 
                 992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b010101; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1211,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b110011; // Expected: {'P': 3213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1212,
                 
                 P
                 , 
                 
                 3213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b111010; // Expected: {'P': 1740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1213,
                 
                 P
                 , 
                 
                 1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b101001; // Expected: {'P': 2173}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1214,
                 
                 P
                 , 
                 
                 2173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100100; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1215,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b101111; // Expected: {'P': 376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1216,
                 
                 P
                 , 
                 
                 376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b111110; // Expected: {'P': 3348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1217,
                 
                 P
                 , 
                 
                 3348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b110011; // Expected: {'P': 1020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1218,
                 
                 P
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b010011; // Expected: {'P': 760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1219,
                 
                 P
                 , 
                 
                 760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b100101; // Expected: {'P': 1036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1220,
                 
                 P
                 , 
                 
                 1036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b101001; // Expected: {'P': 902}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1221,
                 
                 P
                 , 
                 
                 902
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b010011; // Expected: {'P': 323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1222,
                 
                 P
                 , 
                 
                 323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101001; // Expected: {'P': 2378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1223,
                 
                 P
                 , 
                 
                 2378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b000111; // Expected: {'P': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1224,
                 
                 P
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b001011; // Expected: {'P': 594}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1225,
                 
                 P
                 , 
                 
                 594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b111100; // Expected: {'P': 2640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1226,
                 
                 P
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1227,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b110011; // Expected: {'P': 3009}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1228,
                 
                 P
                 , 
                 
                 3009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b111101; // Expected: {'P': 3477}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1229,
                 
                 P
                 , 
                 
                 3477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001011; // Expected: {'P': 374}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1230,
                 
                 P
                 , 
                 
                 374
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100001; // Expected: {'P': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1231,
                 
                 P
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b111110; // Expected: {'P': 248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1232,
                 
                 P
                 , 
                 
                 248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b110110; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1233,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b100100; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1234,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b011000; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1235,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b111000; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1236,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110100; // Expected: {'P': 1664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1237,
                 
                 P
                 , 
                 
                 1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b000110; // Expected: {'P': 312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1238,
                 
                 P
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b111000; // Expected: {'P': 2632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1239,
                 
                 P
                 , 
                 
                 2632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010011; // Expected: {'P': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1240,
                 
                 P
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b011101; // Expected: {'P': 261}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1241,
                 
                 P
                 , 
                 
                 261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b011010; // Expected: {'P': 676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1242,
                 
                 P
                 , 
                 
                 676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b010101; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1243,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100011; // Expected: {'P': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1244,
                 
                 P
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110110; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1245,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b101110; // Expected: {'P': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1246,
                 
                 P
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100011; // Expected: {'P': 1575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1247,
                 
                 P
                 , 
                 
                 1575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b101011; // Expected: {'P': 2451}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1248,
                 
                 P
                 , 
                 
                 2451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1249,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b100101; // Expected: {'P': 2146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1250,
                 
                 P
                 , 
                 
                 2146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b011000; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1251,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b110100; // Expected: {'P': 1300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1252,
                 
                 P
                 , 
                 
                 1300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b010110; // Expected: {'P': 990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1253,
                 
                 P
                 , 
                 
                 990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b100110; // Expected: {'P': 1254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1254,
                 
                 P
                 , 
                 
                 1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b100110; // Expected: {'P': 2128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1255,
                 
                 P
                 , 
                 
                 2128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b100000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1256,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b000010; // Expected: {'P': 14}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1257,
                 
                 P
                 , 
                 
                 14
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b110110; // Expected: {'P': 2484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1258,
                 
                 P
                 , 
                 
                 2484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b110001; // Expected: {'P': 686}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1259,
                 
                 P
                 , 
                 
                 686
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b000001; // Expected: {'P': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1260,
                 
                 P
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b010100; // Expected: {'P': 1040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1261,
                 
                 P
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b101000; // Expected: {'P': 1040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1262,
                 
                 P
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b011101; // Expected: {'P': 348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1263,
                 
                 P
                 , 
                 
                 348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1264,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111001; // Expected: {'P': 2793}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1265,
                 
                 P
                 , 
                 
                 2793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b001111; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1266,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b111100; // Expected: {'P': 3300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1267,
                 
                 P
                 , 
                 
                 3300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b000001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1268,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b101010; // Expected: {'P': 2562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1269,
                 
                 P
                 , 
                 
                 2562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b110011; // Expected: {'P': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1270,
                 
                 P
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100001; // Expected: {'P': 495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1271,
                 
                 P
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b111101; // Expected: {'P': 1342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1272,
                 
                 P
                 , 
                 
                 1342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b110001; // Expected: {'P': 1372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1273,
                 
                 P
                 , 
                 
                 1372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b111110; // Expected: {'P': 1302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1274,
                 
                 P
                 , 
                 
                 1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b000111; // Expected: {'P': 119}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1275,
                 
                 P
                 , 
                 
                 119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b010010; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1276,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b111110; // Expected: {'P': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1277,
                 
                 P
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b011000; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1278,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b001000; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1279,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b110100; // Expected: {'P': 312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1280,
                 
                 P
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b111101; // Expected: {'P': 3294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1281,
                 
                 P
                 , 
                 
                 3294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100000; // Expected: {'P': 1312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1282,
                 
                 P
                 , 
                 
                 1312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b111010; // Expected: {'P': 3596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1283,
                 
                 P
                 , 
                 
                 3596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b001010; // Expected: {'P': 590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1284,
                 
                 P
                 , 
                 
                 590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010001; // Expected: {'P': 952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1285,
                 
                 P
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b010010; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1286,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b001011; // Expected: {'P': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1287,
                 
                 P
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100001; // Expected: {'P': 1353}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1288,
                 
                 P
                 , 
                 
                 1353
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b110111; // Expected: {'P': 2805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1289,
                 
                 P
                 , 
                 
                 2805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b010100; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1290,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b100001; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1291,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b011000; // Expected: {'P': 696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1292,
                 
                 P
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b111001; // Expected: {'P': 342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1293,
                 
                 P
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001001; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1294,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b111010; // Expected: {'P': 1334}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1295,
                 
                 P
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001011; // Expected: {'P': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1296,
                 
                 P
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b111000; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1297,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100010; // Expected: {'P': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1298,
                 
                 P
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b101110; // Expected: {'P': 1058}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1299,
                 
                 P
                 , 
                 
                 1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110011; // Expected: {'P': 153}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1300,
                 
                 P
                 , 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b110110; // Expected: {'P': 2970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1301,
                 
                 P
                 , 
                 
                 2970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b101101; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1302,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010101; // Expected: {'P': 861}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1303,
                 
                 P
                 , 
                 
                 861
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b111010; // Expected: {'P': 580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1304,
                 
                 P
                 , 
                 
                 580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b010001; // Expected: {'P': 476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1305,
                 
                 P
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b001110; // Expected: {'P': 434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1306,
                 
                 P
                 , 
                 
                 434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101110; // Expected: {'P': 1794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1307,
                 
                 P
                 , 
                 
                 1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b101111; // Expected: {'P': 141}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1308,
                 
                 P
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b010011; // Expected: {'P': 494}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1309,
                 
                 P
                 , 
                 
                 494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b000010; // Expected: {'P': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1310,
                 
                 P
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b100001; // Expected: {'P': 396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1311,
                 
                 P
                 , 
                 
                 396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b111011; // Expected: {'P': 3599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1312,
                 
                 P
                 , 
                 
                 3599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011101; // Expected: {'P': 464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1313,
                 
                 P
                 , 
                 
                 464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110111; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1314,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b000101; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1315,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b000111; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1316,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b100010; // Expected: {'P': 2108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1317,
                 
                 P
                 , 
                 
                 2108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001110; // Expected: {'P': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1318,
                 
                 P
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b000110; // Expected: {'P': 102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1319,
                 
                 P
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b011100; // Expected: {'P': 1652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1320,
                 
                 P
                 , 
                 
                 1652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b010000; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1321,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b011111; // Expected: {'P': 1426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1322,
                 
                 P
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b001011; // Expected: {'P': 418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1323,
                 
                 P
                 , 
                 
                 418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b101101; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1324,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b001010; // Expected: {'P': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1325,
                 
                 P
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b110000; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1326,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b100100; // Expected: {'P': 2124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1327,
                 
                 P
                 , 
                 
                 2124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b111010; // Expected: {'P': 290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1328,
                 
                 P
                 , 
                 
                 290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b011000; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1329,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010010; // Expected: {'P': 558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1330,
                 
                 P
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b000011; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1331,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b011110; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1332,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b101110; // Expected: {'P': 1840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1333,
                 
                 P
                 , 
                 
                 1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b011011; // Expected: {'P': 945}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1334,
                 
                 P
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b011101; // Expected: {'P': 1073}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1335,
                 
                 P
                 , 
                 
                 1073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b110101; // Expected: {'P': 1855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1336,
                 
                 P
                 , 
                 
                 1855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100111; // Expected: {'P': 507}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1337,
                 
                 P
                 , 
                 
                 507
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b111110; // Expected: {'P': 1364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1338,
                 
                 P
                 , 
                 
                 1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b001101; // Expected: {'P': 520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1339,
                 
                 P
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100011; // Expected: {'P': 175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1340,
                 
                 P
                 , 
                 
                 175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b111001; // Expected: {'P': 855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1341,
                 
                 P
                 , 
                 
                 855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b000100; // Expected: {'P': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1342,
                 
                 P
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b101111; // Expected: {'P': 2679}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1343,
                 
                 P
                 , 
                 
                 2679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b111000; // Expected: {'P': 3024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1344,
                 
                 P
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b101010; // Expected: {'P': 1386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1345,
                 
                 P
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b000010; // Expected: {'P': 10}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1346,
                 
                 P
                 , 
                 
                 10
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b011010; // Expected: {'P': 1170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1347,
                 
                 P
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b101100; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1348,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b010101; // Expected: {'P': 399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1349,
                 
                 P
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b111101; // Expected: {'P': 3416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1350,
                 
                 P
                 , 
                 
                 3416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b001000; // Expected: {'P': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1351,
                 
                 P
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b011100; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1352,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b010110; // Expected: {'P': 1364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1353,
                 
                 P
                 , 
                 
                 1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b000111; // Expected: {'P': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1354,
                 
                 P
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b000110; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1355,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100101; // Expected: {'P': 1517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1356,
                 
                 P
                 , 
                 
                 1517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b100100; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1357,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b101001; // Expected: {'P': 328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1358,
                 
                 P
                 , 
                 
                 328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b110011; // Expected: {'P': 357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1359,
                 
                 P
                 , 
                 
                 357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b100101; // Expected: {'P': 1258}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1360,
                 
                 P
                 , 
                 
                 1258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1361,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b110111; // Expected: {'P': 2035}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1362,
                 
                 P
                 , 
                 
                 2035
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b011110; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1363,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b000010; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1364,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b001001; // Expected: {'P': 495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1365,
                 
                 P
                 , 
                 
                 495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b101101; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1366,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b101101; // Expected: {'P': 2070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1367,
                 
                 P
                 , 
                 
                 2070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b111011; // Expected: {'P': 1121}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1368,
                 
                 P
                 , 
                 
                 1121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101111; // Expected: {'P': 2350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1369,
                 
                 P
                 , 
                 
                 2350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b011010; // Expected: {'P': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1370,
                 
                 P
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000111; // Expected: {'P': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1371,
                 
                 P
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b111110; // Expected: {'P': 1116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1372,
                 
                 P
                 , 
                 
                 1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b010000; // Expected: {'P': 848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1373,
                 
                 P
                 , 
                 
                 848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b011100; // Expected: {'P': 1372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1374,
                 
                 P
                 , 
                 
                 1372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b110110; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1375,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1376,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b110101; // Expected: {'P': 3233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1377,
                 
                 P
                 , 
                 
                 3233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b111101; // Expected: {'P': 2745}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1378,
                 
                 P
                 , 
                 
                 2745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101100; // Expected: {'P': 2156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1379,
                 
                 P
                 , 
                 
                 2156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000001; // Expected: {'P': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1380,
                 
                 P
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011011; // Expected: {'P': 1377}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1381,
                 
                 P
                 , 
                 
                 1377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b011101; // Expected: {'P': 319}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1382,
                 
                 P
                 , 
                 
                 319
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b110110; // Expected: {'P': 1944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1383,
                 
                 P
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b100111; // Expected: {'P': 546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1384,
                 
                 P
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b001111; // Expected: {'P': 435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1385,
                 
                 P
                 , 
                 
                 435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b111011; // Expected: {'P': 708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1386,
                 
                 P
                 , 
                 
                 708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b000100; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1387,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b101010; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1388,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b100100; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1389,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010000; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1390,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b110101; // Expected: {'P': 265}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1391,
                 
                 P
                 , 
                 
                 265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b110010; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1392,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b011111; // Expected: {'P': 1178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1393,
                 
                 P
                 , 
                 
                 1178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b110010; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1394,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b000111; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1395,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b110111; // Expected: {'P': 1485}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1396,
                 
                 P
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b100110; // Expected: {'P': 1786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1397,
                 
                 P
                 , 
                 
                 1786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101000; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1398,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110011; // Expected: {'P': 2907}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1399,
                 
                 P
                 , 
                 
                 2907
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001100; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1400,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b100010; // Expected: {'P': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1401,
                 
                 P
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b010100; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1402,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b110000; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1403,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b110101; // Expected: {'P': 2915}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1404,
                 
                 P
                 , 
                 
                 2915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000101; // Expected: {'P': 305}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1405,
                 
                 P
                 , 
                 
                 305
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100001; // Expected: {'P': 429}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1406,
                 
                 P
                 , 
                 
                 429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b010011; // Expected: {'P': 722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1407,
                 
                 P
                 , 
                 
                 722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b010010; // Expected: {'P': 666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1408,
                 
                 P
                 , 
                 
                 666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b001111; // Expected: {'P': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1409,
                 
                 P
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b101010; // Expected: {'P': 1974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1410,
                 
                 P
                 , 
                 
                 1974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b111101; // Expected: {'P': 732}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1411,
                 
                 P
                 , 
                 
                 732
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100010; // Expected: {'P': 1394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1412,
                 
                 P
                 , 
                 
                 1394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100000; // Expected: {'P': 864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1413,
                 
                 P
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b111100; // Expected: {'P': 1740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1414,
                 
                 P
                 , 
                 
                 1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b101000; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1415,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b011110; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1416,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b001010; // Expected: {'P': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1417,
                 
                 P
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b001010; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1418,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b011100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1419,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b110110; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1420,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011001; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1421,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b000110; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1422,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111110; // Expected: {'P': 2356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1423,
                 
                 P
                 , 
                 
                 2356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b100010; // Expected: {'P': 544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1424,
                 
                 P
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b000100; // Expected: {'P': 212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1425,
                 
                 P
                 , 
                 
                 212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b000001; // Expected: {'P': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1426,
                 
                 P
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b110111; // Expected: {'P': 1815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1427,
                 
                 P
                 , 
                 
                 1815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b011101; // Expected: {'P': 928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1428,
                 
                 P
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001111; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1429,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b011001; // Expected: {'P': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1430,
                 
                 P
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1431,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010110; // Expected: {'P': 902}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1432,
                 
                 P
                 , 
                 
                 902
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110101; // Expected: {'P': 1643}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1433,
                 
                 P
                 , 
                 
                 1643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1434,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b111001; // Expected: {'P': 2850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1435,
                 
                 P
                 , 
                 
                 2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b101010; // Expected: {'P': 966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1436,
                 
                 P
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b110111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1437,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b011101; // Expected: {'P': 87}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1438,
                 
                 P
                 , 
                 
                 87
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b100111; // Expected: {'P': 117}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1439,
                 
                 P
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b110000; // Expected: {'P': 1728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1440,
                 
                 P
                 , 
                 
                 1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b000101; // Expected: {'P': 55}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1441,
                 
                 P
                 , 
                 
                 55
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b110001; // Expected: {'P': 2205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1442,
                 
                 P
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b001100; // Expected: {'P': 588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1443,
                 
                 P
                 , 
                 
                 588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b000110; // Expected: {'P': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1444,
                 
                 P
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b000100; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1445,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b101000; // Expected: {'P': 1520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1446,
                 
                 P
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111100; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1447,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b000011; // Expected: {'P': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1448,
                 
                 P
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b101111; // Expected: {'P': 2914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1449,
                 
                 P
                 , 
                 
                 2914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b010101; // Expected: {'P': 966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1450,
                 
                 P
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b101000; // Expected: {'P': 2320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1451,
                 
                 P
                 , 
                 
                 2320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b111001; // Expected: {'P': 3534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1452,
                 
                 P
                 , 
                 
                 3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1453,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000011; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1454,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b000001; // Expected: {'P': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1455,
                 
                 P
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b101001; // Expected: {'P': 615}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1456,
                 
                 P
                 , 
                 
                 615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001011; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1457,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b011100; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1458,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110010; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1459,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011111; // Expected: {'P': 1302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1460,
                 
                 P
                 , 
                 
                 1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101000; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1461,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b111000; // Expected: {'P': 3136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1462,
                 
                 P
                 , 
                 
                 3136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b000110; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1463,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101111; // Expected: {'P': 2397}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1464,
                 
                 P
                 , 
                 
                 2397
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b000110; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1465,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b000110; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1466,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b100101; // Expected: {'P': 407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1467,
                 
                 P
                 , 
                 
                 407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b001001; // Expected: {'P': 513}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1468,
                 
                 P
                 , 
                 
                 513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b100000; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1469,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b111001; // Expected: {'P': 1197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1470,
                 
                 P
                 , 
                 
                 1197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b011111; // Expected: {'P': 341}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1471,
                 
                 P
                 , 
                 
                 341
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b101011; // Expected: {'P': 1376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1472,
                 
                 P
                 , 
                 
                 1376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b111101; // Expected: {'P': 2379}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1473,
                 
                 P
                 , 
                 
                 2379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b101101; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1474,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b001000; // Expected: {'P': 320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1475,
                 
                 P
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b100100; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1476,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111011; // Expected: {'P': 2891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1477,
                 
                 P
                 , 
                 
                 2891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b110101; // Expected: {'P': 2597}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1478,
                 
                 P
                 , 
                 
                 2597
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b010100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1479,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b111111; // Expected: {'P': 819}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1480,
                 
                 P
                 , 
                 
                 819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b011000; // Expected: {'P': 312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1481,
                 
                 P
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100000; // Expected: {'P': 416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1482,
                 
                 P
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111001; // Expected: {'P': 3591}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1483,
                 
                 P
                 , 
                 
                 3591
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b001111; // Expected: {'P': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1484,
                 
                 P
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b000110; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1485,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b111111; // Expected: {'P': 1827}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1486,
                 
                 P
                 , 
                 
                 1827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b011000; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1487,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001101; // Expected: {'P': 442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1488,
                 
                 P
                 , 
                 
                 442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b011011; // Expected: {'P': 891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1489,
                 
                 P
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b110110; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1490,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b010011; // Expected: {'P': 1159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1491,
                 
                 P
                 , 
                 
                 1159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b000011; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1492,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100101; // Expected: {'P': 999}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1493,
                 
                 P
                 , 
                 
                 999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1494,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b110110; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1495,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b100000; // Expected: {'P': 1856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1496,
                 
                 P
                 , 
                 
                 1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b010101; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1497,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b001010; // Expected: {'P': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1498,
                 
                 P
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b110101; // Expected: {'P': 636}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1499,
                 
                 P
                 , 
                 
                 636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b110111; // Expected: {'P': 825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1500,
                 
                 P
                 , 
                 
                 825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b010110; // Expected: {'P': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1501,
                 
                 P
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b000011; // Expected: {'P': 42}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1502,
                 
                 P
                 , 
                 
                 42
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b001100; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1503,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b100000; // Expected: {'P': 1024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1504,
                 
                 P
                 , 
                 
                 1024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b001011; // Expected: {'P': 220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1505,
                 
                 P
                 , 
                 
                 220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b010011; // Expected: {'P': 551}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1506,
                 
                 P
                 , 
                 
                 551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b110111; // Expected: {'P': 3410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1507,
                 
                 P
                 , 
                 
                 3410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b101011; // Expected: {'P': 817}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1508,
                 
                 P
                 , 
                 
                 817
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b001001; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1509,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b001000; // Expected: {'P': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1510,
                 
                 P
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b111110; // Expected: {'P': 496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1511,
                 
                 P
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110111; // Expected: {'P': 2145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1512,
                 
                 P
                 , 
                 
                 2145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b001011; // Expected: {'P': 451}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1513,
                 
                 P
                 , 
                 
                 451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b001011; // Expected: {'P': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1514,
                 
                 P
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b011110; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1515,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b101100; // Expected: {'P': 2464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1516,
                 
                 P
                 , 
                 
                 2464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b011011; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1517,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b011000; // Expected: {'P': 1032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1518,
                 
                 P
                 , 
                 
                 1032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b111000; // Expected: {'P': 3192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1519,
                 
                 P
                 , 
                 
                 3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b111110; // Expected: {'P': 868}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1520,
                 
                 P
                 , 
                 
                 868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100000; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1521,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b100111; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1522,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b100000; // Expected: {'P': 1728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1523,
                 
                 P
                 , 
                 
                 1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b111110; // Expected: {'P': 1860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1524,
                 
                 P
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110001; // Expected: {'P': 2646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1525,
                 
                 P
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b111100; // Expected: {'P': 3060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1526,
                 
                 P
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b011100; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1527,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100101; // Expected: {'P': 185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1528,
                 
                 P
                 , 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1529,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b111110; // Expected: {'P': 1488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1530,
                 
                 P
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b111001; // Expected: {'P': 2280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1531,
                 
                 P
                 , 
                 
                 2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b100101; // Expected: {'P': 1628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1532,
                 
                 P
                 , 
                 
                 1628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010010; // Expected: {'P': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1533,
                 
                 P
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b000001; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1534,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b011011; // Expected: {'P': 1053}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1535,
                 
                 P
                 , 
                 
                 1053
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b011000; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1536,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b010100; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1537,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b100010; // Expected: {'P': 1462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1538,
                 
                 P
                 , 
                 
                 1462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b010001; // Expected: {'P': 136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1539,
                 
                 P
                 , 
                 
                 136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b110110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1540,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b101010; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1541,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b001100; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1542,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110111; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1543,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b000011; // Expected: {'P': 138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1544,
                 
                 P
                 , 
                 
                 138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b100111; // Expected: {'P': 1677}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1545,
                 
                 P
                 , 
                 
                 1677
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b100011; // Expected: {'P': 385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1546,
                 
                 P
                 , 
                 
                 385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b011011; // Expected: {'P': 1458}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1547,
                 
                 P
                 , 
                 
                 1458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b011010; // Expected: {'P': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1548,
                 
                 P
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b101010; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1549,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1550,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b001011; // Expected: {'P': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1551,
                 
                 P
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1552,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000011; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1553,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b100111; // Expected: {'P': 1131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1554,
                 
                 P
                 , 
                 
                 1131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b001111; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1555,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b010110; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1556,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b001110; // Expected: {'P': 392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1557,
                 
                 P
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b010000; // Expected: {'P': 368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1558,
                 
                 P
                 , 
                 
                 368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b010001; // Expected: {'P': 255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1559,
                 
                 P
                 , 
                 
                 255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001001; // Expected: {'P': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1560,
                 
                 P
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b000111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1561,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b100111; // Expected: {'P': 2223}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1562,
                 
                 P
                 , 
                 
                 2223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b000010; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1563,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b001100; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1564,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101010; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1565,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b010100; // Expected: {'P': 640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1566,
                 
                 P
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b100011; // Expected: {'P': 1365}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1567,
                 
                 P
                 , 
                 
                 1365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1568,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b001110; // Expected: {'P': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1569,
                 
                 P
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b101010; // Expected: {'P': 2268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1570,
                 
                 P
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b010110; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1571,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b110010; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1572,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b011000; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1573,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110000; // Expected: {'P': 2736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1574,
                 
                 P
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b010011; // Expected: {'P': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1575,
                 
                 P
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b111010; // Expected: {'P': 2552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1576,
                 
                 P
                 , 
                 
                 2552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b100011; // Expected: {'P': 2205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1577,
                 
                 P
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b011001; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1578,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b001001; // Expected: {'P': 9}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1579,
                 
                 P
                 , 
                 
                 9
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b011000; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1580,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b011110; // Expected: {'P': 1770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1581,
                 
                 P
                 , 
                 
                 1770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b101111; // Expected: {'P': 1128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1582,
                 
                 P
                 , 
                 
                 1128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b000111; // Expected: {'P': 441}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1583,
                 
                 P
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b101101; // Expected: {'P': 1845}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1584,
                 
                 P
                 , 
                 
                 1845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100110; // Expected: {'P': 722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1585,
                 
                 P
                 , 
                 
                 722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b001000; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1586,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b101111; // Expected: {'P': 2632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1587,
                 
                 P
                 , 
                 
                 2632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b111010; // Expected: {'P': 2784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1588,
                 
                 P
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b011010; // Expected: {'P': 364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1589,
                 
                 P
                 , 
                 
                 364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b101010; // Expected: {'P': 1050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1590,
                 
                 P
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110111; // Expected: {'P': 3080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1591,
                 
                 P
                 , 
                 
                 3080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b000101; // Expected: {'P': 5}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1592,
                 
                 P
                 , 
                 
                 5
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b100010; // Expected: {'P': 2142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1593,
                 
                 P
                 , 
                 
                 2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b101111; // Expected: {'P': 2115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1594,
                 
                 P
                 , 
                 
                 2115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001111; // Expected: {'P': 345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1595,
                 
                 P
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110010; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1596,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b010000; // Expected: {'P': 832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1597,
                 
                 P
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101000; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1598,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b001111; // Expected: {'P': 855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1599,
                 
                 P
                 , 
                 
                 855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1600,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b101111; // Expected: {'P': 799}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1601,
                 
                 P
                 , 
                 
                 799
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b110101; // Expected: {'P': 1537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1602,
                 
                 P
                 , 
                 
                 1537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100001; // Expected: {'P': 891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1603,
                 
                 P
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b010110; // Expected: {'P': 1100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1604,
                 
                 P
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b011010; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1605,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101010; // Expected: {'P': 2310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1606,
                 
                 P
                 , 
                 
                 2310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b001101; // Expected: {'P': 611}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1607,
                 
                 P
                 , 
                 
                 611
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b011010; // Expected: {'P': 832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1608,
                 
                 P
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001011; // Expected: {'P': 121}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1609,
                 
                 P
                 , 
                 
                 121
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b100101; // Expected: {'P': 2220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1610,
                 
                 P
                 , 
                 
                 2220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b111000; // Expected: {'P': 3304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1611,
                 
                 P
                 , 
                 
                 3304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b010011; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1612,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b001111; // Expected: {'P': 465}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1613,
                 
                 P
                 , 
                 
                 465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110001; // Expected: {'P': 1470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1614,
                 
                 P
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b011011; // Expected: {'P': 486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1615,
                 
                 P
                 , 
                 
                 486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b011000; // Expected: {'P': 1392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1616,
                 
                 P
                 , 
                 
                 1392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110101; // Expected: {'P': 2968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1617,
                 
                 P
                 , 
                 
                 2968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011010; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1618,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b011111; // Expected: {'P': 1395}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1619,
                 
                 P
                 , 
                 
                 1395
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010100; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1620,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b111000; // Expected: {'P': 3248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1621,
                 
                 P
                 , 
                 
                 3248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b101101; // Expected: {'P': 405}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1622,
                 
                 P
                 , 
                 
                 405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b110100; // Expected: {'P': 2392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1623,
                 
                 P
                 , 
                 
                 2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b000001; // Expected: {'P': 35}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1624,
                 
                 P
                 , 
                 
                 35
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100010; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1625,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001101; // Expected: {'P': 650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1626,
                 
                 P
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b011101; // Expected: {'P': 1189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1627,
                 
                 P
                 , 
                 
                 1189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b000101; // Expected: {'P': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1628,
                 
                 P
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b000110; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1629,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b010011; // Expected: {'P': 513}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1630,
                 
                 P
                 , 
                 
                 513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011110; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1631,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b110000; // Expected: {'P': 2784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1632,
                 
                 P
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b101010; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1633,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110010; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1634,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b011111; // Expected: {'P': 1860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1635,
                 
                 P
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b000100; // Expected: {'P': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1636,
                 
                 P
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b101110; // Expected: {'P': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1637,
                 
                 P
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b100110; // Expected: {'P': 304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1638,
                 
                 P
                 , 
                 
                 304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b111101; // Expected: {'P': 3538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1639,
                 
                 P
                 , 
                 
                 3538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001100; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1640,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001110; // Expected: {'P': 602}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1641,
                 
                 P
                 , 
                 
                 602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b011110; // Expected: {'P': 1110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1642,
                 
                 P
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b100010; // Expected: {'P': 1802}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1643,
                 
                 P
                 , 
                 
                 1802
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b100101; // Expected: {'P': 259}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1644,
                 
                 P
                 , 
                 
                 259
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000101; // Expected: {'P': 145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1645,
                 
                 P
                 , 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b010011; // Expected: {'P': 665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1646,
                 
                 P
                 , 
                 
                 665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1647,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b110101; // Expected: {'P': 318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1648,
                 
                 P
                 , 
                 
                 318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101001; // Expected: {'P': 1599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1649,
                 
                 P
                 , 
                 
                 1599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b011101; // Expected: {'P': 1160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1650,
                 
                 P
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b010101; // Expected: {'P': 987}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1651,
                 
                 P
                 , 
                 
                 987
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b011011; // Expected: {'P': 621}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1652,
                 
                 P
                 , 
                 
                 621
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b111000; // Expected: {'P': 1792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1653,
                 
                 P
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b111001; // Expected: {'P': 2565}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1654,
                 
                 P
                 , 
                 
                 2565
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b011100; // Expected: {'P': 1232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1655,
                 
                 P
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100101; // Expected: {'P': 703}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1656,
                 
                 P
                 , 
                 
                 703
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010011; // Expected: {'P': 779}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1657,
                 
                 P
                 , 
                 
                 779
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001000; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1658,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b001001; // Expected: {'P': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1659,
                 
                 P
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b110010; // Expected: {'P': 850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1660,
                 
                 P
                 , 
                 
                 850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b100110; // Expected: {'P': 1292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1661,
                 
                 P
                 , 
                 
                 1292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011011; // Expected: {'P': 648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1662,
                 
                 P
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b100010; // Expected: {'P': 1666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1663,
                 
                 P
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b110010; // Expected: {'P': 1150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1664,
                 
                 P
                 , 
                 
                 1150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b000110; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1665,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b111010; // Expected: {'P': 2900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1666,
                 
                 P
                 , 
                 
                 2900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b010100; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1667,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b001101; // Expected: {'P': 546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1668,
                 
                 P
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b011101; // Expected: {'P': 406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1669,
                 
                 P
                 , 
                 
                 406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b110011; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1670,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b100010; // Expected: {'P': 102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1671,
                 
                 P
                 , 
                 
                 102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b010010; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1672,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101111; // Expected: {'P': 2961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1673,
                 
                 P
                 , 
                 
                 2961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010001; // Expected: {'P': 527}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1674,
                 
                 P
                 , 
                 
                 527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101001; // Expected: {'P': 2255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1675,
                 
                 P
                 , 
                 
                 2255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b111001; // Expected: {'P': 1767}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1676,
                 
                 P
                 , 
                 
                 1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1677,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101110; // Expected: {'P': 506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1678,
                 
                 P
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010100; // Expected: {'P': 820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1679,
                 
                 P
                 , 
                 
                 820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b000111; // Expected: {'P': 273}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1680,
                 
                 P
                 , 
                 
                 273
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b111110; // Expected: {'P': 1240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1681,
                 
                 P
                 , 
                 
                 1240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b011011; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1682,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b100111; // Expected: {'P': 819}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1683,
                 
                 P
                 , 
                 
                 819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b001110; // Expected: {'P': 490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1684,
                 
                 P
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b011110; // Expected: {'P': 1050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1685,
                 
                 P
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b000101; // Expected: {'P': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1686,
                 
                 P
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111101; // Expected: {'P': 976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1687,
                 
                 P
                 , 
                 
                 976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b010101; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1688,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b001100; // Expected: {'P': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1689,
                 
                 P
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001000; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1690,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b111111; // Expected: {'P': 945}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1691,
                 
                 P
                 , 
                 
                 945
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b100001; // Expected: {'P': 825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1692,
                 
                 P
                 , 
                 
                 825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b100000; // Expected: {'P': 928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1693,
                 
                 P
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b001010; // Expected: {'P': 520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1694,
                 
                 P
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000111; // Expected: {'P': 266}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1695,
                 
                 P
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111000; // Expected: {'P': 2744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1696,
                 
                 P
                 , 
                 
                 2744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b010110; // Expected: {'P': 1122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1697,
                 
                 P
                 , 
                 
                 1122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b010111; // Expected: {'P': 1426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1698,
                 
                 P
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b111100; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1699,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b010111; // Expected: {'P': 874}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1700,
                 
                 P
                 , 
                 
                 874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100011; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1701,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111010; // Expected: {'P': 3654}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1702,
                 
                 P
                 , 
                 
                 3654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b110101; // Expected: {'P': 1802}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1703,
                 
                 P
                 , 
                 
                 1802
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b111000; // Expected: {'P': 392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1704,
                 
                 P
                 , 
                 
                 392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b001011; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1705,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b011011; // Expected: {'P': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1706,
                 
                 P
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b011010; // Expected: {'P': 1144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1707,
                 
                 P
                 , 
                 
                 1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110111; // Expected: {'P': 2915}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1708,
                 
                 P
                 , 
                 
                 2915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b111000; // Expected: {'P': 1232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1709,
                 
                 P
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b111101; // Expected: {'P': 1464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1710,
                 
                 P
                 , 
                 
                 1464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b100110; // Expected: {'P': 912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1711,
                 
                 P
                 , 
                 
                 912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b001101; // Expected: {'P': 130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1712,
                 
                 P
                 , 
                 
                 130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b001101; // Expected: {'P': 507}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1713,
                 
                 P
                 , 
                 
                 507
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b010110; // Expected: {'P': 352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1714,
                 
                 P
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b011000; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1715,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b011001; // Expected: {'P': 1500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1716,
                 
                 P
                 , 
                 
                 1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001010; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1717,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b010010; // Expected: {'P': 414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1718,
                 
                 P
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111111; // Expected: {'P': 2646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1719,
                 
                 P
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b101111; // Expected: {'P': 2820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1720,
                 
                 P
                 , 
                 
                 2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b110110; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1721,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100011; // Expected: {'P': 1470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1722,
                 
                 P
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b111010; // Expected: {'P': 812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1723,
                 
                 P
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011011; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1724,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110011; // Expected: {'P': 510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1725,
                 
                 P
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b001111; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1726,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b001110; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1727,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111011; // Expected: {'P': 2242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1728,
                 
                 P
                 , 
                 
                 2242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b011000; // Expected: {'P': 1104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1729,
                 
                 P
                 , 
                 
                 1104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b011000; // Expected: {'P': 1272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1730,
                 
                 P
                 , 
                 
                 1272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001010; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1731,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b111010; // Expected: {'P': 928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1732,
                 
                 P
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1733,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b101010; // Expected: {'P': 1554}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1734,
                 
                 P
                 , 
                 
                 1554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b001001; // Expected: {'P': 459}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1735,
                 
                 P
                 , 
                 
                 459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b111010; // Expected: {'P': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1736,
                 
                 P
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b101111; // Expected: {'P': 658}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1737,
                 
                 P
                 , 
                 
                 658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b110100; // Expected: {'P': 2132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1738,
                 
                 P
                 , 
                 
                 2132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100001; // Expected: {'P': 1518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1739,
                 
                 P
                 , 
                 
                 1518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b001010; // Expected: {'P': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1740,
                 
                 P
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b010100; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1741,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b010110; // Expected: {'P': 506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1742,
                 
                 P
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b110011; // Expected: {'P': 969}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1743,
                 
                 P
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b001000; // Expected: {'P': 312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1744,
                 
                 P
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110000; // Expected: {'P': 2544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1745,
                 
                 P
                 , 
                 
                 2544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b001101; // Expected: {'P': 741}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1746,
                 
                 P
                 , 
                 
                 741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b001000; // Expected: {'P': 456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1747,
                 
                 P
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b010110; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1748,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111111; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1749,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b000001; // Expected: {'P': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 1750,
                 
                 P
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b111100; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1751,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b101010; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1752,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b101011; // Expected: {'P': 215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1753,
                 
                 P
                 , 
                 
                 215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b010101; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1754,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b010111; // Expected: {'P': 184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1755,
                 
                 P
                 , 
                 
                 184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b111001; // Expected: {'P': 1938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1756,
                 
                 P
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b011010; // Expected: {'P': 754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1757,
                 
                 P
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111010; // Expected: {'P': 2204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1758,
                 
                 P
                 , 
                 
                 2204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b101110; // Expected: {'P': 2208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1759,
                 
                 P
                 , 
                 
                 2208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011000; // Expected: {'P': 1224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1760,
                 
                 P
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b001001; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1761,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b101100; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1762,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b011100; // Expected: {'P': 476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1763,
                 
                 P
                 , 
                 
                 476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b011011; // Expected: {'P': 783}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1764,
                 
                 P
                 , 
                 
                 783
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b101010; // Expected: {'P': 2604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1765,
                 
                 P
                 , 
                 
                 2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b001000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1766,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b011010; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1767,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b111000; // Expected: {'P': 1960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1768,
                 
                 P
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b001000; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1769,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1770,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b000111; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1771,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b010011; // Expected: {'P': 1026}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1772,
                 
                 P
                 , 
                 
                 1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b111011; // Expected: {'P': 2773}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1773,
                 
                 P
                 , 
                 
                 2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b011100; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1774,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b101110; // Expected: {'P': 1150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1775,
                 
                 P
                 , 
                 
                 1150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b011110; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1776,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b100110; // Expected: {'P': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1777,
                 
                 P
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b111111; // Expected: {'P': 2709}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1778,
                 
                 P
                 , 
                 
                 2709
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b011010; // Expected: {'P': 988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1779,
                 
                 P
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b000010; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1780,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b100011; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1781,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001000; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1782,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b101001; // Expected: {'P': 1517}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1783,
                 
                 P
                 , 
                 
                 1517
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b111000; // Expected: {'P': 1064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1784,
                 
                 P
                 , 
                 
                 1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b010110; // Expected: {'P': 814}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1785,
                 
                 P
                 , 
                 
                 814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b001011; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1786,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b011011; // Expected: {'P': 1485}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1787,
                 
                 P
                 , 
                 
                 1485
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b100111; // Expected: {'P': 1560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1788,
                 
                 P
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001101; // Expected: {'P': 793}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 1789,
                 
                 P
                 , 
                 
                 793
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b101101; // Expected: {'P': 1350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1790,
                 
                 P
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b110011; // Expected: {'P': 663}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1791,
                 
                 P
                 , 
                 
                 663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b101001; // Expected: {'P': 1025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1792,
                 
                 P
                 , 
                 
                 1025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b001010; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1793,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b011000; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1794,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b101001; // Expected: {'P': 2296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1795,
                 
                 P
                 , 
                 
                 2296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110100; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1796,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1797,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b011010; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1798,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b010110; // Expected: {'P': 374}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1799,
                 
                 P
                 , 
                 
                 374
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b000101; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1800,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b000101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1801,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b100011; // Expected: {'P': 525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1802,
                 
                 P
                 , 
                 
                 525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b010010; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1803,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b100101; // Expected: {'P': 629}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1804,
                 
                 P
                 , 
                 
                 629
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1805,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b100101; // Expected: {'P': 740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1806,
                 
                 P
                 , 
                 
                 740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b010110; // Expected: {'P': 1254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1807,
                 
                 P
                 , 
                 
                 1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b010111; // Expected: {'P': 322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1808,
                 
                 P
                 , 
                 
                 322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b101100; // Expected: {'P': 2376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1809,
                 
                 P
                 , 
                 
                 2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b011111; // Expected: {'P': 558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1810,
                 
                 P
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b010001; // Expected: {'P': 680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1811,
                 
                 P
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b101000; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1812,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b100110; // Expected: {'P': 76}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1813,
                 
                 P
                 , 
                 
                 76
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b110001; // Expected: {'P': 2548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1814,
                 
                 P
                 , 
                 
                 2548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b100101; // Expected: {'P': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1815,
                 
                 P
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b101010; // Expected: {'P': 1344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1816,
                 
                 P
                 , 
                 
                 1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b100101; // Expected: {'P': 2294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1817,
                 
                 P
                 , 
                 
                 2294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b001100; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1818,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b010011; // Expected: {'P': 475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1819,
                 
                 P
                 , 
                 
                 475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b100111; // Expected: {'P': 2106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1820,
                 
                 P
                 , 
                 
                 2106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b001010; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1821,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b001011; // Expected: {'P': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1822,
                 
                 P
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001010; // Expected: {'P': 610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1823,
                 
                 P
                 , 
                 
                 610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b010001; // Expected: {'P': 816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1824,
                 
                 P
                 , 
                 
                 816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b111000; // Expected: {'P': 1904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1825,
                 
                 P
                 , 
                 
                 1904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b101010; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1826,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b000011; // Expected: {'P': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1827,
                 
                 P
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b010110; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1828,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b111011; // Expected: {'P': 3068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 1829,
                 
                 P
                 , 
                 
                 3068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b010010; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1830,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b100010; // Expected: {'P': 2006}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1831,
                 
                 P
                 , 
                 
                 2006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110100; // Expected: {'P': 2756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1832,
                 
                 P
                 , 
                 
                 2756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b100000; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1833,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b001111; // Expected: {'P': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1834,
                 
                 P
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b100011; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1835,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b011111; // Expected: {'P': 1674}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1836,
                 
                 P
                 , 
                 
                 1674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b011010; // Expected: {'P': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1837,
                 
                 P
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b001111; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1838,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b001100; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1839,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b011001; // Expected: {'P': 325}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1840,
                 
                 P
                 , 
                 
                 325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100110; // Expected: {'P': 1748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1841,
                 
                 P
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b111010; // Expected: {'P': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1842,
                 
                 P
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b110010; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1843,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b111001; // Expected: {'P': 1653}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1844,
                 
                 P
                 , 
                 
                 1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b100101; // Expected: {'P': 1776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1845,
                 
                 P
                 , 
                 
                 1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b011101; // Expected: {'P': 580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1846,
                 
                 P
                 , 
                 
                 580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b111101; // Expected: {'P': 122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 1847,
                 
                 P
                 , 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b011010; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1848,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b001001; // Expected: {'P': 297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1849,
                 
                 P
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000100; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1850,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b101000; // Expected: {'P': 1000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1851,
                 
                 P
                 , 
                 
                 1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b001001; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1852,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b000111; // Expected: {'P': 203}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1853,
                 
                 P
                 , 
                 
                 203
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b101110; // Expected: {'P': 2484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 1854,
                 
                 P
                 , 
                 
                 2484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b101000; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1855,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b000110; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1856,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b110111; // Expected: {'P': 1210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1857,
                 
                 P
                 , 
                 
                 1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b100000; // Expected: {'P': 256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1858,
                 
                 P
                 , 
                 
                 256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b010111; // Expected: {'P': 897}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1859,
                 
                 P
                 , 
                 
                 897
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b101101; // Expected: {'P': 2790}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1860,
                 
                 P
                 , 
                 
                 2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001010; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1861,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b011000; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1862,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b000010; // Expected: {'P': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1863,
                 
                 P
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b011110; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1864,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b110100; // Expected: {'P': 1144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1865,
                 
                 P
                 , 
                 
                 1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b101010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 1866,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b011011; // Expected: {'P': 1161}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1867,
                 
                 P
                 , 
                 
                 1161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001001; // Expected: {'P': 207}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1868,
                 
                 P
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b001111; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1869,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b011010; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1870,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b010001; // Expected: {'P': 17}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1871,
                 
                 P
                 , 
                 
                 17
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b010100; // Expected: {'P': 680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1872,
                 
                 P
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b000111; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1873,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010011; // Expected: {'P': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1874,
                 
                 P
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b011100; // Expected: {'P': 532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1875,
                 
                 P
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b011001; // Expected: {'P': 1225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1876,
                 
                 P
                 , 
                 
                 1225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110110; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 1877,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011011; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1878,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b111110; // Expected: {'P': 1550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1879,
                 
                 P
                 , 
                 
                 1550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100100; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1880,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110100; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 1881,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b010111; // Expected: {'P': 782}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1882,
                 
                 P
                 , 
                 
                 782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b000100; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1883,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b110111; // Expected: {'P': 990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1884,
                 
                 P
                 , 
                 
                 990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b010101; // Expected: {'P': 1113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1885,
                 
                 P
                 , 
                 
                 1113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b111001; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1886,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b001100; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1887,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b100000; // Expected: {'P': 1376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1888,
                 
                 P
                 , 
                 
                 1376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b110001; // Expected: {'P': 1715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1889,
                 
                 P
                 , 
                 
                 1715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b111110; // Expected: {'P': 310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1890,
                 
                 P
                 , 
                 
                 310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011000; // Expected: {'P': 1128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 1891,
                 
                 P
                 , 
                 
                 1128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b001110; // Expected: {'P': 364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1892,
                 
                 P
                 , 
                 
                 364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110000; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1893,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b010100; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1894,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b101111; // Expected: {'P': 1927}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1895,
                 
                 P
                 , 
                 
                 1927
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b011100; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1896,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110111; // Expected: {'P': 1705}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1897,
                 
                 P
                 , 
                 
                 1705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b010100; // Expected: {'P': 740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 1898,
                 
                 P
                 , 
                 
                 740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b010111; // Expected: {'P': 851}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1899,
                 
                 P
                 , 
                 
                 851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b100010; // Expected: {'P': 952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1900,
                 
                 P
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b000100; // Expected: {'P': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 1901,
                 
                 P
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b111110; // Expected: {'P': 2232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 1902,
                 
                 P
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b011010; // Expected: {'P': 884}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1903,
                 
                 P
                 , 
                 
                 884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b000101; // Expected: {'P': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1904,
                 
                 P
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b000101; // Expected: {'P': 285}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1905,
                 
                 P
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b100101; // Expected: {'P': 925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 1906,
                 
                 P
                 , 
                 
                 925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b101000; // Expected: {'P': 1880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1907,
                 
                 P
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b010001; // Expected: {'P': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1908,
                 
                 P
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b010101; // Expected: {'P': 294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1909,
                 
                 P
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b100010; // Expected: {'P': 1768}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1910,
                 
                 P
                 , 
                 
                 1768
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b011110; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 1911,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b001100; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1912,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111010; // Expected: {'P': 2842}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 1913,
                 
                 P
                 , 
                 
                 2842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b010000; // Expected: {'P': 352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1914,
                 
                 P
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110111; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 1915,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b001011; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1916,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b010010; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1917,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b010110; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1918,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b001010; // Expected: {'P': 550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1919,
                 
                 P
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110010; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 1920,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010101; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 1921,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b111001; // Expected: {'P': 114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1922,
                 
                 P
                 , 
                 
                 114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001011; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 1923,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000110; // Expected: {'P': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1924,
                 
                 P
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b101001; // Expected: {'P': 738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1925,
                 
                 P
                 , 
                 
                 738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010011; // Expected: {'P': 1064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 1926,
                 
                 P
                 , 
                 
                 1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b100000; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 1927,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b110011; // Expected: {'P': 612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1928,
                 
                 P
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b011010; // Expected: {'P': 1534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1929,
                 
                 P
                 , 
                 
                 1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b100011; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 1930,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b001001; // Expected: {'P': 369}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1931,
                 
                 P
                 , 
                 
                 369
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b011010; // Expected: {'P': 1066}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 1932,
                 
                 P
                 , 
                 
                 1066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b110101; // Expected: {'P': 901}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 1933,
                 
                 P
                 , 
                 
                 901
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b000110; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1934,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b010010; // Expected: {'P': 1062}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 1935,
                 
                 P
                 , 
                 
                 1062
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b000010; // Expected: {'P': 28}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1936,
                 
                 P
                 , 
                 
                 28
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000110; // Expected: {'P': 366}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1937,
                 
                 P
                 , 
                 
                 366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b101000; // Expected: {'P': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1938,
                 
                 P
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b010000; // Expected: {'P': 944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1939,
                 
                 P
                 , 
                 
                 944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101001; // Expected: {'P': 2050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 1940,
                 
                 P
                 , 
                 
                 2050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b011111; // Expected: {'P': 62}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1941,
                 
                 P
                 , 
                 
                 62
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b000111; // Expected: {'P': 301}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1942,
                 
                 P
                 , 
                 
                 301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b000010; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1943,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b100111; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1944,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b000110; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1945,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b001010; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 1946,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b010000; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 1947,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001110; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1948,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b000101; // Expected: {'P': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 1949,
                 
                 P
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1950,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b001111; // Expected: {'P': 75}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 1951,
                 
                 P
                 , 
                 
                 75
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b011101; // Expected: {'P': 1711}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1952,
                 
                 P
                 , 
                 
                 1711
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b111001; // Expected: {'P': 2052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1953,
                 
                 P
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b000111; // Expected: {'P': 77}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1954,
                 
                 P
                 , 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b101000; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 1955,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b100111; // Expected: {'P': 702}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1956,
                 
                 P
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b101100; // Expected: {'P': 2024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 1957,
                 
                 P
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b111111; // Expected: {'P': 1701}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1958,
                 
                 P
                 , 
                 
                 1701
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b101101; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1959,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b101011; // Expected: {'P': 1548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 1960,
                 
                 P
                 , 
                 
                 1548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b001110; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 1961,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001100; // Expected: {'P': 276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 1962,
                 
                 P
                 , 
                 
                 276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b001001; // Expected: {'P': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1963,
                 
                 P
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100111; // Expected: {'P': 1755}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1964,
                 
                 P
                 , 
                 
                 1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100100; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 1965,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b001001; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 1966,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b000011; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 1967,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101111; // Expected: {'P': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 1968,
                 
                 P
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b111000; // Expected: {'P': 784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 1969,
                 
                 P
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b111100; // Expected: {'P': 2400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1970,
                 
                 P
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b001000; // Expected: {'P': 256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 1971,
                 
                 P
                 , 
                 
                 256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1972,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111111; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 1973,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b110011; // Expected: {'P': 2295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 1974,
                 
                 P
                 , 
                 
                 2295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b011111; // Expected: {'P': 713}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 1975,
                 
                 P
                 , 
                 
                 713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b100010; // Expected: {'P': 1938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 1976,
                 
                 P
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b110000; // Expected: {'P': 1776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 1977,
                 
                 P
                 , 
                 
                 1776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b111100; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1978,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b011101; // Expected: {'P': 1334}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1979,
                 
                 P
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b100110; // Expected: {'P': 874}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 1980,
                 
                 P
                 , 
                 
                 874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b011100; // Expected: {'P': 644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 1981,
                 
                 P
                 , 
                 
                 644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b000110; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 1982,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b010001; // Expected: {'P': 1020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 1983,
                 
                 P
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b000111; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 1984,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b101101; // Expected: {'P': 810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 1985,
                 
                 P
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b100001; // Expected: {'P': 1287}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1986,
                 
                 P
                 , 
                 
                 1287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000010; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 1987,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b010110; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 1988,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b111001; // Expected: {'P': 1425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 1989,
                 
                 P
                 , 
                 
                 1425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b011011; // Expected: {'P': 1647}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 1990,
                 
                 P
                 , 
                 
                 1647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b110001; // Expected: {'P': 3038}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 1991,
                 
                 P
                 , 
                 
                 3038
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 1992,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b100001; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 1993,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b111100; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1994,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111100; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 1995,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b011001; // Expected: {'P': 1125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 1996,
                 
                 P
                 , 
                 
                 1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b100111; // Expected: {'P': 741}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 1997,
                 
                 P
                 , 
                 
                 741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b011101; // Expected: {'P': 522}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 1998,
                 
                 P
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b010111; // Expected: {'P': 667}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 1999,
                 
                 P
                 , 
                 
                 667
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011101; // Expected: {'P': 1363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2000,
                 
                 P
                 , 
                 
                 1363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b010110; // Expected: {'P': 638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2001,
                 
                 P
                 , 
                 
                 638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b101001; // Expected: {'P': 1968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2002,
                 
                 P
                 , 
                 
                 1968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b111000; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2003,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2004,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b111111; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2005,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111001; // Expected: {'P': 2622}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 2006,
                 
                 P
                 , 
                 
                 2622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b010101; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2007,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110101; // Expected: {'P': 477}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2008,
                 
                 P
                 , 
                 
                 477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110101; // Expected: {'P': 2067}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2009,
                 
                 P
                 , 
                 
                 2067
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b000001; // Expected: {'P': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2010,
                 
                 P
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b001011; // Expected: {'P': 693}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2011,
                 
                 P
                 , 
                 
                 693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b101001; // Expected: {'P': 1927}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2012,
                 
                 P
                 , 
                 
                 1927
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b001111; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2013,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b000101; // Expected: {'P': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2014,
                 
                 P
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b111111; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2015,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b110001; // Expected: {'P': 1764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2016,
                 
                 P
                 , 
                 
                 1764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b110000; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2017,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b010010; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2018,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b101100; // Expected: {'P': 1100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2019,
                 
                 P
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b010011; // Expected: {'P': 1197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2020,
                 
                 P
                 , 
                 
                 1197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b101110; // Expected: {'P': 1012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2021,
                 
                 P
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b100110; // Expected: {'P': 1938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2022,
                 
                 P
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b000101; // Expected: {'P': 185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2023,
                 
                 P
                 , 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b001000; // Expected: {'P': 496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2024,
                 
                 P
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b001111; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2025,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100001; // Expected: {'P': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2026,
                 
                 P
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b001010; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 2027,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b100001; // Expected: {'P': 1881}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2028,
                 
                 P
                 , 
                 
                 1881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b001111; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2029,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b110000; // Expected: {'P': 2832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2030,
                 
                 P
                 , 
                 
                 2832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b011011; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2031,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b110000; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2032,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b110011; // Expected: {'P': 3060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2033,
                 
                 P
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010000; // Expected: {'P': 656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2034,
                 
                 P
                 , 
                 
                 656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b010011; // Expected: {'P': 646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2035,
                 
                 P
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b111010; // Expected: {'P': 1276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2036,
                 
                 P
                 , 
                 
                 1276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b001111; // Expected: {'P': 405}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2037,
                 
                 P
                 , 
                 
                 405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b011110; // Expected: {'P': 1470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2038,
                 
                 P
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b111001; // Expected: {'P': 1311}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 2039,
                 
                 P
                 , 
                 
                 1311
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b001111; // Expected: {'P': 810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2040,
                 
                 P
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b111110; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2041,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b111010; // Expected: {'P': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2042,
                 
                 P
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b000101; // Expected: {'P': 205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2043,
                 
                 P
                 , 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b000101; // Expected: {'P': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2044,
                 
                 P
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b010111; // Expected: {'P': 1357}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2045,
                 
                 P
                 , 
                 
                 1357
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b010111; // Expected: {'P': 920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2046,
                 
                 P
                 , 
                 
                 920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b011001; // Expected: {'P': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 2047,
                 
                 P
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b111011; // Expected: {'P': 2183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2048,
                 
                 P
                 , 
                 
                 2183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b011011; // Expected: {'P': 837}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2049,
                 
                 P
                 , 
                 
                 837
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b010011; // Expected: {'P': 285}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2050,
                 
                 P
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b110111; // Expected: {'P': 1925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2051,
                 
                 P
                 , 
                 
                 1925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011100; // Expected: {'P': 448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2052,
                 
                 P
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b101110; // Expected: {'P': 690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2053,
                 
                 P
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b000011; // Expected: {'P': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2054,
                 
                 P
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b110001; // Expected: {'P': 980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2055,
                 
                 P
                 , 
                 
                 980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b000101; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2056,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b011100; // Expected: {'P': 1568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2057,
                 
                 P
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b010011; // Expected: {'P': 817}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2058,
                 
                 P
                 , 
                 
                 817
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b101011; // Expected: {'P': 1634}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2059,
                 
                 P
                 , 
                 
                 1634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011000; // Expected: {'P': 576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2060,
                 
                 P
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b101010; // Expected: {'P': 1848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2061,
                 
                 P
                 , 
                 
                 1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b001001; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2062,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b000111; // Expected: {'P': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 2063,
                 
                 P
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b010000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2064,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b100111; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2065,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b000101; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2066,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000010; // Expected: {'P': 16}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2067,
                 
                 P
                 , 
                 
                 16
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b010111; // Expected: {'P': 1104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2068,
                 
                 P
                 , 
                 
                 1104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110110; // Expected: {'P': 486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2069,
                 
                 P
                 , 
                 
                 486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b100001; // Expected: {'P': 1782}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2070,
                 
                 P
                 , 
                 
                 1782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b100001; // Expected: {'P': 363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2071,
                 
                 P
                 , 
                 
                 363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b100111; // Expected: {'P': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2072,
                 
                 P
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b111010; // Expected: {'P': 2320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2073,
                 
                 P
                 , 
                 
                 2320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b001101; // Expected: {'P': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2074,
                 
                 P
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b010111; // Expected: {'P': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2075,
                 
                 P
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b111110; // Expected: {'P': 1612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2076,
                 
                 P
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000100; // Expected: {'P': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2077,
                 
                 P
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b100011; // Expected: {'P': 980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2078,
                 
                 P
                 , 
                 
                 980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111101; // Expected: {'P': 2562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2079,
                 
                 P
                 , 
                 
                 2562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2080,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b001001; // Expected: {'P': 171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2081,
                 
                 P
                 , 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b111101; // Expected: {'P': 1037}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2082,
                 
                 P
                 , 
                 
                 1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b101001; // Expected: {'P': 984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2083,
                 
                 P
                 , 
                 
                 984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100111; // Expected: {'P': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2084,
                 
                 P
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010000; // Expected: {'P': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2085,
                 
                 P
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b010100; // Expected: {'P': 420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2086,
                 
                 P
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b111110; // Expected: {'P': 3100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2087,
                 
                 P
                 , 
                 
                 3100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b111101; // Expected: {'P': 1281}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2088,
                 
                 P
                 , 
                 
                 1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110101; // Expected: {'P': 3021}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2089,
                 
                 P
                 , 
                 
                 3021
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b001110; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2090,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b111010; // Expected: {'P': 2146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2091,
                 
                 P
                 , 
                 
                 2146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b101101; // Expected: {'P': 765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 2092,
                 
                 P
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b011110; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2093,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b110011; // Expected: {'P': 1377}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2094,
                 
                 P
                 , 
                 
                 1377
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b001110; // Expected: {'P': 448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2095,
                 
                 P
                 , 
                 
                 448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101110; // Expected: {'P': 322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2096,
                 
                 P
                 , 
                 
                 322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b001011; // Expected: {'P': 396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2097,
                 
                 P
                 , 
                 
                 396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b001100; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2098,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b001110; // Expected: {'P': 588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2099,
                 
                 P
                 , 
                 
                 588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100100; // Expected: {'P': 1620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2100,
                 
                 P
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101111; // Expected: {'P': 47}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2101,
                 
                 P
                 , 
                 
                 47
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b101000; // Expected: {'P': 1240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2102,
                 
                 P
                 , 
                 
                 1240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b101011; // Expected: {'P': 2623}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2103,
                 
                 P
                 , 
                 
                 2623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100000; // Expected: {'P': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2104,
                 
                 P
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b100100; // Expected: {'P': 1296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2105,
                 
                 P
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b101110; // Expected: {'P': 598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2106,
                 
                 P
                 , 
                 
                 598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b111000; // Expected: {'P': 1736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2107,
                 
                 P
                 , 
                 
                 1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b001100; // Expected: {'P': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2108,
                 
                 P
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2109,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010100; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2110,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b010000; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2111,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011000; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2112,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b101100; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2113,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b011101; // Expected: {'P': 1537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2114,
                 
                 P
                 , 
                 
                 1537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b100000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2115,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b010001; // Expected: {'P': 85}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2116,
                 
                 P
                 , 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b010001; // Expected: {'P': 1003}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2117,
                 
                 P
                 , 
                 
                 1003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b000111; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 2118,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110011; // Expected: {'P': 1224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2119,
                 
                 P
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b110001; // Expected: {'P': 2107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2120,
                 
                 P
                 , 
                 
                 2107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101101; // Expected: {'P': 1575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 2121,
                 
                 P
                 , 
                 
                 1575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b001111; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2122,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110001; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2123,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b000001; // Expected: {'P': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2124,
                 
                 P
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b011100; // Expected: {'P': 1596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2125,
                 
                 P
                 , 
                 
                 1596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b110110; // Expected: {'P': 2754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2126,
                 
                 P
                 , 
                 
                 2754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b101010; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2127,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b110110; // Expected: {'P': 2322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2128,
                 
                 P
                 , 
                 
                 2322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000011; // Expected: {'P': 177}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2129,
                 
                 P
                 , 
                 
                 177
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b000011; // Expected: {'P': 141}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2130,
                 
                 P
                 , 
                 
                 141
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010001; // Expected: {'P': 748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2131,
                 
                 P
                 , 
                 
                 748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b110111; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2132,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b110101; // Expected: {'P': 2544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2133,
                 
                 P
                 , 
                 
                 2544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b100000; // Expected: {'P': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2134,
                 
                 P
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b111110; // Expected: {'P': 3038}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2135,
                 
                 P
                 , 
                 
                 3038
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b010001; // Expected: {'P': 697}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2136,
                 
                 P
                 , 
                 
                 697
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b101100; // Expected: {'P': 792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2137,
                 
                 P
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2138,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b100000; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2139,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b111000; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2140,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101110; // Expected: {'P': 2392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2141,
                 
                 P
                 , 
                 
                 2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b000100; // Expected: {'P': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2142,
                 
                 P
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101111; // Expected: {'P': 752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2143,
                 
                 P
                 , 
                 
                 752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b011101; // Expected: {'P': 145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2144,
                 
                 P
                 , 
                 
                 145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b010010; // Expected: {'P': 936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2145,
                 
                 P
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b101001; // Expected: {'P': 1189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2146,
                 
                 P
                 , 
                 
                 1189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b000101; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2147,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111001; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 2148,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b000110; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2149,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111101; // Expected: {'P': 549}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2150,
                 
                 P
                 , 
                 
                 549
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b110010; // Expected: {'P': 1900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2151,
                 
                 P
                 , 
                 
                 1900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b100111; // Expected: {'P': 2457}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2152,
                 
                 P
                 , 
                 
                 2457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b100000; // Expected: {'P': 1280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2153,
                 
                 P
                 , 
                 
                 1280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b101011; // Expected: {'P': 1591}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2154,
                 
                 P
                 , 
                 
                 1591
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b000010; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2155,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b111100; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2156,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b110010; // Expected: {'P': 1100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2157,
                 
                 P
                 , 
                 
                 1100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b110111; // Expected: {'P': 1870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2158,
                 
                 P
                 , 
                 
                 1870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000011; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2159,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b001000; // Expected: {'P': 376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2160,
                 
                 P
                 , 
                 
                 376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011010; // Expected: {'P': 1222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2161,
                 
                 P
                 , 
                 
                 1222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b010100; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2162,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111101; // Expected: {'P': 3843}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2163,
                 
                 P
                 , 
                 
                 3843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b000010; // Expected: {'P': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2164,
                 
                 P
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2165,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111100; // Expected: {'P': 3600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2166,
                 
                 P
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b000011; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2167,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b001101; // Expected: {'P': 780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2168,
                 
                 P
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b101001; // Expected: {'P': 943}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2169,
                 
                 P
                 , 
                 
                 943
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110010; // Expected: {'P': 1500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2170,
                 
                 P
                 , 
                 
                 1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b111011; // Expected: {'P': 2301}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2171,
                 
                 P
                 , 
                 
                 2301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b011111; // Expected: {'P': 1240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2172,
                 
                 P
                 , 
                 
                 1240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010011; // Expected: {'P': 133}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2173,
                 
                 P
                 , 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b110000; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2174,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b100110; // Expected: {'P': 1558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2175,
                 
                 P
                 , 
                 
                 1558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b111100; // Expected: {'P': 3240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2176,
                 
                 P
                 , 
                 
                 3240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b111000; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2177,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001000; // Expected: {'P': 272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2178,
                 
                 P
                 , 
                 
                 272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b010111; // Expected: {'P': 1380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2179,
                 
                 P
                 , 
                 
                 1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b111110; // Expected: {'P': 620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2180,
                 
                 P
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b101100; // Expected: {'P': 1716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2181,
                 
                 P
                 , 
                 
                 1716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b011111; // Expected: {'P': 1736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2182,
                 
                 P
                 , 
                 
                 1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b110000; // Expected: {'P': 2304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2183,
                 
                 P
                 , 
                 
                 2304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b000010; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2184,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b111011; // Expected: {'P': 2832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2185,
                 
                 P
                 , 
                 
                 2832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b001000; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2186,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b100101; // Expected: {'P': 444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2187,
                 
                 P
                 , 
                 
                 444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b000011; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2188,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b010011; // Expected: {'P': 437}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2189,
                 
                 P
                 , 
                 
                 437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b011111; // Expected: {'P': 496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2190,
                 
                 P
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b001101; // Expected: {'P': 403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2191,
                 
                 P
                 , 
                 
                 403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b001000; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2192,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b100101; // Expected: {'P': 1480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2193,
                 
                 P
                 , 
                 
                 1480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001001; // Expected: {'P': 549}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2194,
                 
                 P
                 , 
                 
                 549
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b011011; // Expected: {'P': 1701}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2195,
                 
                 P
                 , 
                 
                 1701
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2196,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b100100; // Expected: {'P': 1368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2197,
                 
                 P
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b010110; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2198,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001001; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2199,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b000101; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2200,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b010111; // Expected: {'P': 1311}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2201,
                 
                 P
                 , 
                 
                 1311
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b100101; // Expected: {'P': 962}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2202,
                 
                 P
                 , 
                 
                 962
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b010110; // Expected: {'P': 770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2203,
                 
                 P
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b001101; // Expected: {'P': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2204,
                 
                 P
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b111111; // Expected: {'P': 1449}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2205,
                 
                 P
                 , 
                 
                 1449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b101101; // Expected: {'P': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 2206,
                 
                 P
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b100000; // Expected: {'P': 992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2207,
                 
                 P
                 , 
                 
                 992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100011; // Expected: {'P': 1610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2208,
                 
                 P
                 , 
                 
                 1610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b100010; // Expected: {'P': 34}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 2209,
                 
                 P
                 , 
                 
                 34
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b111100; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2210,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b011000; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2211,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b001111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2212,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b001110; // Expected: {'P': 322}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2213,
                 
                 P
                 , 
                 
                 322
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b101101; // Expected: {'P': 855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 2214,
                 
                 P
                 , 
                 
                 855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b110101; // Expected: {'P': 2332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2215,
                 
                 P
                 , 
                 
                 2332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001101; // Expected: {'P': 208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2216,
                 
                 P
                 , 
                 
                 208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b110011; // Expected: {'P': 2958}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2217,
                 
                 P
                 , 
                 
                 2958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b011110; // Expected: {'P': 990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2218,
                 
                 P
                 , 
                 
                 990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b111001; // Expected: {'P': 570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 2219,
                 
                 P
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b110101; // Expected: {'P': 2014}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2220,
                 
                 P
                 , 
                 
                 2014
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b010111; // Expected: {'P': 1035}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2221,
                 
                 P
                 , 
                 
                 1035
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b011110; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2222,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b101111; // Expected: {'P': 2021}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2223,
                 
                 P
                 , 
                 
                 2021
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b010110; // Expected: {'P': 1210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2224,
                 
                 P
                 , 
                 
                 1210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b100100; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2225,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b000011; // Expected: {'P': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2226,
                 
                 P
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b010111; // Expected: {'P': 1334}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2227,
                 
                 P
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b010111; // Expected: {'P': 1403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2228,
                 
                 P
                 , 
                 
                 1403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b100011; // Expected: {'P': 1785}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2229,
                 
                 P
                 , 
                 
                 1785
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b101100; // Expected: {'P': 2596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2230,
                 
                 P
                 , 
                 
                 2596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b011110; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2231,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b000001; // Expected: {'P': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2232,
                 
                 P
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000011; // Expected: {'P': 183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2233,
                 
                 P
                 , 
                 
                 183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b010000; // Expected: {'P': 736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2234,
                 
                 P
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b011001; // Expected: {'P': 975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 2235,
                 
                 P
                 , 
                 
                 975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2236,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b110000; // Expected: {'P': 2352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2237,
                 
                 P
                 , 
                 
                 2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b111100; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2238,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b001110; // Expected: {'P': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2239,
                 
                 P
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b101100; // Expected: {'P': 396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2240,
                 
                 P
                 , 
                 
                 396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b101011; // Expected: {'P': 2365}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2241,
                 
                 P
                 , 
                 
                 2365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b110100; // Expected: {'P': 2444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2242,
                 
                 P
                 , 
                 
                 2444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b011100; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2243,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110100; // Expected: {'P': 1612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2244,
                 
                 P
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b110110; // Expected: {'P': 1620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2245,
                 
                 P
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b100100; // Expected: {'P': 1692}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2246,
                 
                 P
                 , 
                 
                 1692
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b100110; // Expected: {'P': 608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2247,
                 
                 P
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b101001; // Expected: {'P': 205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2248,
                 
                 P
                 , 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b111010; // Expected: {'P': 986}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2249,
                 
                 P
                 , 
                 
                 986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b001100; // Expected: {'P': 492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2250,
                 
                 P
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b011111; // Expected: {'P': 744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2251,
                 
                 P
                 , 
                 
                 744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b001001; // Expected: {'P': 558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2252,
                 
                 P
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b010101; // Expected: {'P': 1281}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2253,
                 
                 P
                 , 
                 
                 1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101111; // Expected: {'P': 2444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2254,
                 
                 P
                 , 
                 
                 2444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b100100; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2255,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b001111; // Expected: {'P': 780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2256,
                 
                 P
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b111111; // Expected: {'P': 2961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2257,
                 
                 P
                 , 
                 
                 2961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b100000; // Expected: {'P': 1216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2258,
                 
                 P
                 , 
                 
                 1216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b110001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2259,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b100111; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2260,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b101100; // Expected: {'P': 1628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2261,
                 
                 P
                 , 
                 
                 1628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b011111; // Expected: {'P': 992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2262,
                 
                 P
                 , 
                 
                 992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b101101; // Expected: {'P': 585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 2263,
                 
                 P
                 , 
                 
                 585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b011100; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2264,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000010; // Expected: {'P': 122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2265,
                 
                 P
                 , 
                 
                 122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b001001; // Expected: {'P': 261}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2266,
                 
                 P
                 , 
                 
                 261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b001110; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2267,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100101; // Expected: {'P': 1554}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2268,
                 
                 P
                 , 
                 
                 1554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b011110; // Expected: {'P': 1140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2269,
                 
                 P
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b110010; // Expected: {'P': 650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2270,
                 
                 P
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b101011; // Expected: {'P': 1118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2271,
                 
                 P
                 , 
                 
                 1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110010; // Expected: {'P': 1550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2272,
                 
                 P
                 , 
                 
                 1550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111110; // Expected: {'P': 3720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2273,
                 
                 P
                 , 
                 
                 3720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b000111; // Expected: {'P': 329}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 2274,
                 
                 P
                 , 
                 
                 329
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b001000; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2275,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100001; // Expected: {'P': 1221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2276,
                 
                 P
                 , 
                 
                 1221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b101111; // Expected: {'P': 2538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2277,
                 
                 P
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b101010; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2278,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b110100; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2279,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b010000; // Expected: {'P': 608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2280,
                 
                 P
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b000010; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2281,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100100; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2282,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b111100; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2283,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b111110; // Expected: {'P': 1922}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2284,
                 
                 P
                 , 
                 
                 1922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b000001; // Expected: {'P': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2285,
                 
                 P
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b000110; // Expected: {'P': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2286,
                 
                 P
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b010011; // Expected: {'P': 1083}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2287,
                 
                 P
                 , 
                 
                 1083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b010001; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2288,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100110; // Expected: {'P': 1710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2289,
                 
                 P
                 , 
                 
                 1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b001100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2290,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b100111; // Expected: {'P': 1521}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2291,
                 
                 P
                 , 
                 
                 1521
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b110000; // Expected: {'P': 912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2292,
                 
                 P
                 , 
                 
                 912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b010000; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2293,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101010; // Expected: {'P': 2142}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2294,
                 
                 P
                 , 
                 
                 2142
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b110011; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2295,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b110010; // Expected: {'P': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2296,
                 
                 P
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b011111; // Expected: {'P': 1054}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2297,
                 
                 P
                 , 
                 
                 1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b111010; // Expected: {'P': 2668}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2298,
                 
                 P
                 , 
                 
                 2668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b010010; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2299,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b101100; // Expected: {'P': 2684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2300,
                 
                 P
                 , 
                 
                 2684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b001001; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2301,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b100111; // Expected: {'P': 1053}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2302,
                 
                 P
                 , 
                 
                 1053
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010110; // Expected: {'P': 286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2303,
                 
                 P
                 , 
                 
                 286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b101111; // Expected: {'P': 1269}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2304,
                 
                 P
                 , 
                 
                 1269
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b110101; // Expected: {'P': 2491}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2305,
                 
                 P
                 , 
                 
                 2491
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2306,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b111111; // Expected: {'P': 1638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2307,
                 
                 P
                 , 
                 
                 1638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b010101; // Expected: {'P': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2308,
                 
                 P
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b101100; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2309,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b111000; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2310,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b110110; // Expected: {'P': 2106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2311,
                 
                 P
                 , 
                 
                 2106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b101001; // Expected: {'P': 410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2312,
                 
                 P
                 , 
                 
                 410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b001011; // Expected: {'P': 506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2313,
                 
                 P
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b001011; // Expected: {'P': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2314,
                 
                 P
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b100101; // Expected: {'P': 2072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2315,
                 
                 P
                 , 
                 
                 2072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b010111; // Expected: {'P': 1196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2316,
                 
                 P
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b110110; // Expected: {'P': 1242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2317,
                 
                 P
                 , 
                 
                 1242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b001011; // Expected: {'P': 275}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2318,
                 
                 P
                 , 
                 
                 275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b000011; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2319,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b000011; // Expected: {'P': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2320,
                 
                 P
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101000; // Expected: {'P': 2080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2321,
                 
                 P
                 , 
                 
                 2080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101011; // Expected: {'P': 1505}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2322,
                 
                 P
                 , 
                 
                 1505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b010101; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2323,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b100111; // Expected: {'P': 2262}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2324,
                 
                 P
                 , 
                 
                 2262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b010111; // Expected: {'P': 276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2325,
                 
                 P
                 , 
                 
                 276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b101000; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2326,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b010011; // Expected: {'P': 684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2327,
                 
                 P
                 , 
                 
                 684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b011011; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2328,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b101100; // Expected: {'P': 2288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2329,
                 
                 P
                 , 
                 
                 2288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b101100; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2330,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b001100; // Expected: {'P': 516}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2331,
                 
                 P
                 , 
                 
                 516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b110111; // Expected: {'P': 550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2332,
                 
                 P
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b010110; // Expected: {'P': 1386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2333,
                 
                 P
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b001101; // Expected: {'P': 728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2334,
                 
                 P
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b001110; // Expected: {'P': 658}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2335,
                 
                 P
                 , 
                 
                 658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b001001; // Expected: {'P': 477}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2336,
                 
                 P
                 , 
                 
                 477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b101100; // Expected: {'P': 1540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2337,
                 
                 P
                 , 
                 
                 1540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b011011; // Expected: {'P': 1539}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2338,
                 
                 P
                 , 
                 
                 1539
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b010111; // Expected: {'P': 690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2339,
                 
                 P
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b001011; // Expected: {'P': 605}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2340,
                 
                 P
                 , 
                 
                 605
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b111011; // Expected: {'P': 1062}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2341,
                 
                 P
                 , 
                 
                 1062
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b011000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2342,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110001; // Expected: {'P': 441}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2343,
                 
                 P
                 , 
                 
                 441
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111110; // Expected: {'P': 558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2344,
                 
                 P
                 , 
                 
                 558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b111100; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2345,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b011101; // Expected: {'P': 1624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2346,
                 
                 P
                 , 
                 
                 1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b101010; // Expected: {'P': 1428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2347,
                 
                 P
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000110; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2348,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b011101; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2349,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b100111; // Expected: {'P': 663}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2350,
                 
                 P
                 , 
                 
                 663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b001100; // Expected: {'P': 240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2351,
                 
                 P
                 , 
                 
                 240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b110100; // Expected: {'P': 728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2352,
                 
                 P
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b111111; // Expected: {'P': 2016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2353,
                 
                 P
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b111101; // Expected: {'P': 2318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2354,
                 
                 P
                 , 
                 
                 2318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b110001; // Expected: {'P': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2355,
                 
                 P
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2356,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b010111; // Expected: {'P': 1288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2357,
                 
                 P
                 , 
                 
                 1288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b000010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2358,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b001000; // Expected: {'P': 416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2359,
                 
                 P
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101000; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2360,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b000111; // Expected: {'P': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 2361,
                 
                 P
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b100100; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2362,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b000010; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2363,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b011111; // Expected: {'P': 1922}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2364,
                 
                 P
                 , 
                 
                 1922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b101111; // Expected: {'P': 893}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2365,
                 
                 P
                 , 
                 
                 893
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b101111; // Expected: {'P': 2773}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2366,
                 
                 P
                 , 
                 
                 2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b001101; // Expected: {'P': 91}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2367,
                 
                 P
                 , 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b110100; // Expected: {'P': 3120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2368,
                 
                 P
                 , 
                 
                 3120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b011111; // Expected: {'P': 1457}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2369,
                 
                 P
                 , 
                 
                 1457
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b111011; // Expected: {'P': 3658}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2370,
                 
                 P
                 , 
                 
                 3658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b010110; // Expected: {'P': 594}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2371,
                 
                 P
                 , 
                 
                 594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b101110; // Expected: {'P': 782}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2372,
                 
                 P
                 , 
                 
                 782
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b100001; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2373,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b110110; // Expected: {'P': 2646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2374,
                 
                 P
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b001100; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2375,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b110110; // Expected: {'P': 864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2376,
                 
                 P
                 , 
                 
                 864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b110111; // Expected: {'P': 2640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2377,
                 
                 P
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b110010; // Expected: {'P': 1450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2378,
                 
                 P
                 , 
                 
                 1450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b100000; // Expected: {'P': 1344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2379,
                 
                 P
                 , 
                 
                 1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b001101; // Expected: {'P': 494}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2380,
                 
                 P
                 , 
                 
                 494
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b100011; // Expected: {'P': 2135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2381,
                 
                 P
                 , 
                 
                 2135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b010111; // Expected: {'P': 299}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2382,
                 
                 P
                 , 
                 
                 299
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100110; // Expected: {'P': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2383,
                 
                 P
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b010011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2384,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b110101; // Expected: {'P': 848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2385,
                 
                 P
                 , 
                 
                 848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b110001; // Expected: {'P': 1519}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2386,
                 
                 P
                 , 
                 
                 1519
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b101100; // Expected: {'P': 1672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2387,
                 
                 P
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b000100; // Expected: {'P': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2388,
                 
                 P
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b101001; // Expected: {'P': 1558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2389,
                 
                 P
                 , 
                 
                 1558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b011010; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2390,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b010100; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2391,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b101000; // Expected: {'P': 640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2392,
                 
                 P
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b011100; // Expected: {'P': 728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2393,
                 
                 P
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b011101; // Expected: {'P': 957}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2394,
                 
                 P
                 , 
                 
                 957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100011; // Expected: {'P': 455}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2395,
                 
                 P
                 , 
                 
                 455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110010; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2396,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b000110; // Expected: {'P': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2397,
                 
                 P
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b001000; // Expected: {'P': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2398,
                 
                 P
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b100100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2399,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b110011; // Expected: {'P': 561}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2400,
                 
                 P
                 , 
                 
                 561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b101011; // Expected: {'P': 559}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2401,
                 
                 P
                 , 
                 
                 559
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b011110; // Expected: {'P': 1170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2402,
                 
                 P
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b110000; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2403,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b010110; // Expected: {'P': 198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2404,
                 
                 P
                 , 
                 
                 198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b011111; // Expected: {'P': 1581}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2405,
                 
                 P
                 , 
                 
                 1581
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010111; // Expected: {'P': 713}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2406,
                 
                 P
                 , 
                 
                 713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b111000; // Expected: {'P': 1848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2407,
                 
                 P
                 , 
                 
                 1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b101001; // Expected: {'P': 1107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2408,
                 
                 P
                 , 
                 
                 1107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b011011; // Expected: {'P': 27}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2409,
                 
                 P
                 , 
                 
                 27
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b001110; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2410,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b111100; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2411,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b010100; // Expected: {'P': 200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2412,
                 
                 P
                 , 
                 
                 200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b101100; // Expected: {'P': 1804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2413,
                 
                 P
                 , 
                 
                 1804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2414,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b011111; // Expected: {'P': 1023}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2415,
                 
                 P
                 , 
                 
                 1023
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010000; B = 6'b100001; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010000; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2416,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b000110; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2417,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b101011; // Expected: {'P': 2107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2418,
                 
                 P
                 , 
                 
                 2107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b100110; // Expected: {'P': 988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2419,
                 
                 P
                 , 
                 
                 988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b111010; // Expected: {'P': 1102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2420,
                 
                 P
                 , 
                 
                 1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b000110; // Expected: {'P': 30}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2421,
                 
                 P
                 , 
                 
                 30
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b001110; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2422,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b111010; // Expected: {'P': 1160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2423,
                 
                 P
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b111110; // Expected: {'P': 1736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2424,
                 
                 P
                 , 
                 
                 1736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001101; // Expected: {'P': 143}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2425,
                 
                 P
                 , 
                 
                 143
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010100; // Expected: {'P': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2426,
                 
                 P
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b010000; // Expected: {'P': 752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2427,
                 
                 P
                 , 
                 
                 752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b010100; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2428,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b101000; // Expected: {'P': 1160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2429,
                 
                 P
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b100100; // Expected: {'P': 1836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2430,
                 
                 P
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b100101; // Expected: {'P': 1665}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2431,
                 
                 P
                 , 
                 
                 1665
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b100101; // Expected: {'P': 666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2432,
                 
                 P
                 , 
                 
                 666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b100110; // Expected: {'P': 2280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2433,
                 
                 P
                 , 
                 
                 2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b011110; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2434,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101010; // Expected: {'P': 2646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2435,
                 
                 P
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b010101; // Expected: {'P': 567}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2436,
                 
                 P
                 , 
                 
                 567
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b101110; // Expected: {'P': 2300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2437,
                 
                 P
                 , 
                 
                 2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b100111; // Expected: {'P': 1170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2438,
                 
                 P
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b111111; // Expected: {'P': 2331}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b111111; | Outputs: P=%b | Expected: P=%d",
                 2439,
                 
                 P
                 , 
                 
                 2331
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2440,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b011101; // Expected: {'P': 1450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2441,
                 
                 P
                 , 
                 
                 1450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2442,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b010110; // Expected: {'P': 1034}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2443,
                 
                 P
                 , 
                 
                 1034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b101000; // Expected: {'P': 1640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b101000; | Outputs: P=%b | Expected: P=%d",
                 2444,
                 
                 P
                 , 
                 
                 1640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b110010; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2445,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b110101; // Expected: {'P': 2703}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2446,
                 
                 P
                 , 
                 
                 2703
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b001111; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2447,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111011; // Expected: {'P': 2478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2448,
                 
                 P
                 , 
                 
                 2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b010001; // Expected: {'P': 986}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2449,
                 
                 P
                 , 
                 
                 986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101001; // Expected: {'P': 2583}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2450,
                 
                 P
                 , 
                 
                 2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2451,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b101001; // Expected: {'P': 2091}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2452,
                 
                 P
                 , 
                 
                 2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b110110; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b110110; | Outputs: P=%b | Expected: P=%d",
                 2453,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b101010; // Expected: {'P': 1302}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b101010; | Outputs: P=%b | Expected: P=%d",
                 2454,
                 
                 P
                 , 
                 
                 1302
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110010; B = 6'b110111; // Expected: {'P': 2750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2455,
                 
                 P
                 , 
                 
                 2750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b110101; // Expected: {'P': 2756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2456,
                 
                 P
                 , 
                 
                 2756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b001010; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 2457,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b011100; // Expected: {'P': 224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2458,
                 
                 P
                 , 
                 
                 224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b010100; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2459,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110011; B = 6'b001000; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110011; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2460,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b010101; // Expected: {'P': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2461,
                 
                 P
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b000011; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2462,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b001101; // Expected: {'P': 169}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2463,
                 
                 P
                 , 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b000100; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2464,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b011011; // Expected: {'P': 1296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2465,
                 
                 P
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110000; // Expected: {'P': 432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2466,
                 
                 P
                 , 
                 
                 432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b001101; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2467,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110011; // Expected: {'P': 1632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2468,
                 
                 P
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b000101; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2469,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b011111; // Expected: {'P': 837}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2470,
                 
                 P
                 , 
                 
                 837
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010000; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2471,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010111; B = 6'b010101; // Expected: {'P': 483}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010111; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2472,
                 
                 P
                 , 
                 
                 483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b011100; // Expected: {'P': 1036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2473,
                 
                 P
                 , 
                 
                 1036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b011000; // Expected: {'P': 984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2474,
                 
                 P
                 , 
                 
                 984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b111101; // Expected: {'P': 2257}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2475,
                 
                 P
                 , 
                 
                 2257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b011000; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2476,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b110000; // Expected: {'P': 2256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2477,
                 
                 P
                 , 
                 
                 2256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b010011; // Expected: {'P': 627}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2478,
                 
                 P
                 , 
                 
                 627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110111; // Expected: {'P': 2970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2479,
                 
                 P
                 , 
                 
                 2970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b111010; // Expected: {'P': 1218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2480,
                 
                 P
                 , 
                 
                 1218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b101011; // Expected: {'P': 1419}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2481,
                 
                 P
                 , 
                 
                 1419
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b010001; // Expected: {'P': 595}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2482,
                 
                 P
                 , 
                 
                 595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100111; B = 6'b000011; // Expected: {'P': 117}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100111; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2483,
                 
                 P
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b010010; // Expected: {'P': 576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2484,
                 
                 P
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100111; // Expected: {'P': 1794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2485,
                 
                 P
                 , 
                 
                 1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b100000; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2486,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b101100; // Expected: {'P': 968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2487,
                 
                 P
                 , 
                 
                 968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b000101; // Expected: {'P': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2488,
                 
                 P
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b100110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2489,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b001000; // Expected: {'P': 424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2490,
                 
                 P
                 , 
                 
                 424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011101; B = 6'b010010; // Expected: {'P': 522}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011101; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2491,
                 
                 P
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b100100; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2492,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b100110; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2493,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b110101; // Expected: {'P': 1272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2494,
                 
                 P
                 , 
                 
                 1272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000100; B = 6'b101011; // Expected: {'P': 172}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000100; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2495,
                 
                 P
                 , 
                 
                 172
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b000001; // Expected: {'P': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2496,
                 
                 P
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2497,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b100001; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2498,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b100010; // Expected: {'P': 1904}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 2499,
                 
                 P
                 , 
                 
                 1904
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000101; B = 6'b010110; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000101; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2500,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b101011; // Expected: {'P': 860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2501,
                 
                 P
                 , 
                 
                 860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b110010; // Expected: {'P': 2850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2502,
                 
                 P
                 , 
                 
                 2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b001011; // Expected: {'P': 187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2503,
                 
                 P
                 , 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001111; // Expected: {'P': 915}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2504,
                 
                 P
                 , 
                 
                 915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b001101; // Expected: {'P': 39}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2505,
                 
                 P
                 , 
                 
                 39
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100011; // Expected: {'P': 1295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2506,
                 
                 P
                 , 
                 
                 1295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b010110; // Expected: {'P': 682}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2507,
                 
                 P
                 , 
                 
                 682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b110101; // Expected: {'P': 53}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2508,
                 
                 P
                 , 
                 
                 53
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101111; B = 6'b000100; // Expected: {'P': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101111; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2509,
                 
                 P
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b111001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 2510,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b100011; // Expected: {'P': 2065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2511,
                 
                 P
                 , 
                 
                 2065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110010; // Expected: {'P': 2700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2512,
                 
                 P
                 , 
                 
                 2700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b100001; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2513,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b101111; // Expected: {'P': 987}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b101111; | Outputs: P=%b | Expected: P=%d",
                 2514,
                 
                 P
                 , 
                 
                 987
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b100001; // Expected: {'P': 1254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2515,
                 
                 P
                 , 
                 
                 1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b101101; // Expected: {'P': 2025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b101101; | Outputs: P=%b | Expected: P=%d",
                 2516,
                 
                 P
                 , 
                 
                 2025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010101; // Expected: {'P': 147}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2517,
                 
                 P
                 , 
                 
                 147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b110011; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2518,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b111101; // Expected: {'P': 2196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2519,
                 
                 P
                 , 
                 
                 2196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b011111; // Expected: {'P': 1519}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2520,
                 
                 P
                 , 
                 
                 1519
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b101110; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2521,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b100001; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b100001; | Outputs: P=%b | Expected: P=%d",
                 2522,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b000010; // Expected: {'P': 74}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2523,
                 
                 P
                 , 
                 
                 74
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101000; B = 6'b111000; // Expected: {'P': 2240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101000; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2524,
                 
                 P
                 , 
                 
                 2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b111011; // Expected: {'P': 3540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2525,
                 
                 P
                 , 
                 
                 3540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b011101; // Expected: {'P': 725}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2526,
                 
                 P
                 , 
                 
                 725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b011011; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2527,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b010100; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2528,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b110101; // Expected: {'P': 424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2529,
                 
                 P
                 , 
                 
                 424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b000100; // Expected: {'P': 148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2530,
                 
                 P
                 , 
                 
                 148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b111110; // Expected: {'P': 3224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2531,
                 
                 P
                 , 
                 
                 3224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b110101; // Expected: {'P': 1378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2532,
                 
                 P
                 , 
                 
                 1378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b001111; // Expected: {'P': 930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2533,
                 
                 P
                 , 
                 
                 930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b110101; // Expected: {'P': 2809}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2534,
                 
                 P
                 , 
                 
                 2809
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b111100; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b111100; | Outputs: P=%b | Expected: P=%d",
                 2535,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b011111; // Expected: {'P': 465}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2536,
                 
                 P
                 , 
                 
                 465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b111110; // Expected: {'P': 2294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2537,
                 
                 P
                 , 
                 
                 2294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b110001; // Expected: {'P': 1029}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b110001; | Outputs: P=%b | Expected: P=%d",
                 2538,
                 
                 P
                 , 
                 
                 1029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b010010; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2539,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b011100; // Expected: {'P': 1484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b011100; | Outputs: P=%b | Expected: P=%d",
                 2540,
                 
                 P
                 , 
                 
                 1484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b010001; // Expected: {'P': 1037}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2541,
                 
                 P
                 , 
                 
                 1037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001011; B = 6'b001111; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001011; B = 6'b001111; | Outputs: P=%b | Expected: P=%d",
                 2542,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b010000; // Expected: {'P': 416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2543,
                 
                 P
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b001010; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b001010; | Outputs: P=%b | Expected: P=%d",
                 2544,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b101100; // Expected: {'P': 1364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2545,
                 
                 P
                 , 
                 
                 1364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b001110; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2546,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b010000; // Expected: {'P': 976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b010000; | Outputs: P=%b | Expected: P=%d",
                 2547,
                 
                 P
                 , 
                 
                 976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000111; B = 6'b010111; // Expected: {'P': 161}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000111; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2548,
                 
                 P
                 , 
                 
                 161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b110101; // Expected: {'P': 1113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2549,
                 
                 P
                 , 
                 
                 1113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b011010; // Expected: {'P': 1612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2550,
                 
                 P
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2551,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110000; B = 6'b011010; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110000; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2552,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001001; B = 6'b110011; // Expected: {'P': 459}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001001; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2553,
                 
                 P
                 , 
                 
                 459
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b001110; // Expected: {'P': 196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2554,
                 
                 P
                 , 
                 
                 196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b001110; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2555,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b100000; // Expected: {'P': 1888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2556,
                 
                 P
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b110010; // Expected: {'P': 2450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2557,
                 
                 P
                 , 
                 
                 2450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011001; B = 6'b010001; // Expected: {'P': 425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011001; B = 6'b010001; | Outputs: P=%b | Expected: P=%d",
                 2558,
                 
                 P
                 , 
                 
                 425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b001000; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2559,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b000110; // Expected: {'P': 276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2560,
                 
                 P
                 , 
                 
                 276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b110010; // Expected: {'P': 2950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2561,
                 
                 P
                 , 
                 
                 2950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2562,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b001000; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b001000; | Outputs: P=%b | Expected: P=%d",
                 2563,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b010101; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2564,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b110010; // Expected: {'P': 2250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2565,
                 
                 P
                 , 
                 
                 2250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011100; B = 6'b011001; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011100; B = 6'b011001; | Outputs: P=%b | Expected: P=%d",
                 2566,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b000111; // Expected: {'P': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b000111; | Outputs: P=%b | Expected: P=%d",
                 2567,
                 
                 P
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b101100; // Expected: {'P': 1936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b101100; | Outputs: P=%b | Expected: P=%d",
                 2568,
                 
                 P
                 , 
                 
                 1936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b110111; // Expected: {'P': 3190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b110111; | Outputs: P=%b | Expected: P=%d",
                 2569,
                 
                 P
                 , 
                 
                 3190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b110011; // Expected: {'P': 1683}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b110011; | Outputs: P=%b | Expected: P=%d",
                 2570,
                 
                 P
                 , 
                 
                 1683
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b111110; // Expected: {'P': 930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2571,
                 
                 P
                 , 
                 
                 930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001101; B = 6'b100010; // Expected: {'P': 442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001101; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 2572,
                 
                 P
                 , 
                 
                 442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b000011; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2573,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b000100; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2574,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b001110; // Expected: {'P': 644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2575,
                 
                 P
                 , 
                 
                 644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111010; B = 6'b000100; // Expected: {'P': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111010; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2576,
                 
                 P
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b001101; // Expected: {'P': 195}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2577,
                 
                 P
                 , 
                 
                 195
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b000010; // Expected: {'P': 92}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2578,
                 
                 P
                 , 
                 
                 92
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b110100; // Expected: {'P': 2548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2579,
                 
                 P
                 , 
                 
                 2548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b111010; // Expected: {'P': 2436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2580,
                 
                 P
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b101001; // Expected: {'P': 1763}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b101001; | Outputs: P=%b | Expected: P=%d",
                 2581,
                 
                 P
                 , 
                 
                 1763
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b111011; // Expected: {'P': 3304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2582,
                 
                 P
                 , 
                 
                 3304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101001; B = 6'b111011; // Expected: {'P': 2419}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101001; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2583,
                 
                 P
                 , 
                 
                 2419
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001111; B = 6'b001001; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001111; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2584,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b100110; // Expected: {'P': 2242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2585,
                 
                 P
                 , 
                 
                 2242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b111011; // Expected: {'P': 354}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2586,
                 
                 P
                 , 
                 
                 354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011000; B = 6'b000100; // Expected: {'P': 96}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011000; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2587,
                 
                 P
                 , 
                 
                 96
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110001; B = 6'b011010; // Expected: {'P': 1274}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110001; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2588,
                 
                 P
                 , 
                 
                 1274
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001000; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001000; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2589,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001110; B = 6'b101110; // Expected: {'P': 644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001110; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2590,
                 
                 P
                 , 
                 
                 644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b000110; // Expected: {'P': 318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2591,
                 
                 P
                 , 
                 
                 318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b100011; // Expected: {'P': 1155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2592,
                 
                 P
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110111; B = 6'b111011; // Expected: {'P': 3245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110111; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2593,
                 
                 P
                 , 
                 
                 3245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b101110; // Expected: {'P': 2898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b101110; | Outputs: P=%b | Expected: P=%d",
                 2594,
                 
                 P
                 , 
                 
                 2898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b011101; // Expected: {'P': 290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b011101; | Outputs: P=%b | Expected: P=%d",
                 2595,
                 
                 P
                 , 
                 
                 290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010101; B = 6'b100011; // Expected: {'P': 735}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010101; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2596,
                 
                 P
                 , 
                 
                 735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b111001; // Expected: {'P': 3021}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b111001; | Outputs: P=%b | Expected: P=%d",
                 2597,
                 
                 P
                 , 
                 
                 3021
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001100; B = 6'b100110; // Expected: {'P': 456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001100; B = 6'b100110; | Outputs: P=%b | Expected: P=%d",
                 2598,
                 
                 P
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b000001; // Expected: {'P': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2599,
                 
                 P
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100011; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100011; | Outputs: P=%b | Expected: P=%d",
                 2600,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111110; B = 6'b000101; // Expected: {'P': 310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111110; B = 6'b000101; | Outputs: P=%b | Expected: P=%d",
                 2601,
                 
                 P
                 , 
                 
                 310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111111; B = 6'b111110; // Expected: {'P': 3906}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111111; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2602,
                 
                 P
                 , 
                 
                 3906
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b001100; // Expected: {'P': 732}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2603,
                 
                 P
                 , 
                 
                 732
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011111; B = 6'b100111; // Expected: {'P': 1209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011111; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2604,
                 
                 P
                 , 
                 
                 1209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b001101; // Expected: {'P': 585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b001101; | Outputs: P=%b | Expected: P=%d",
                 2605,
                 
                 P
                 , 
                 
                 585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100011; B = 6'b100101; // Expected: {'P': 1295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2606,
                 
                 P
                 , 
                 
                 1295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010011; B = 6'b000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010011; B = 6'b000000; | Outputs: P=%b | Expected: P=%d",
                 2607,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b001100; // Expected: {'P': 312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2608,
                 
                 P
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b010010; // Expected: {'P': 1026}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2609,
                 
                 P
                 , 
                 
                 1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b001110; // Expected: {'P': 532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2610,
                 
                 P
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011110; B = 6'b100000; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2611,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b011000; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b011000; | Outputs: P=%b | Expected: P=%d",
                 2612,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000001; B = 6'b000010; // Expected: {'P': 2}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000001; B = 6'b000010; | Outputs: P=%b | Expected: P=%d",
                 2613,
                 
                 P
                 , 
                 
                 2
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b001001; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b001001; | Outputs: P=%b | Expected: P=%d",
                 2614,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b011010; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2615,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100100; B = 6'b011111; // Expected: {'P': 1116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100100; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2616,
                 
                 P
                 , 
                 
                 1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b111010; // Expected: {'P': 3132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2617,
                 
                 P
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011010; B = 6'b000110; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011010; B = 6'b000110; | Outputs: P=%b | Expected: P=%d",
                 2618,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b111000; // Expected: {'P': 2464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b111000; | Outputs: P=%b | Expected: P=%d",
                 2619,
                 
                 P
                 , 
                 
                 2464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110100; B = 6'b110010; // Expected: {'P': 2600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110100; B = 6'b110010; | Outputs: P=%b | Expected: P=%d",
                 2620,
                 
                 P
                 , 
                 
                 2600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b001110; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b001110; | Outputs: P=%b | Expected: P=%d",
                 2621,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b110100; // Expected: {'P': 1040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2622,
                 
                 P
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b111101; // Expected: {'P': 366}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b111101; | Outputs: P=%b | Expected: P=%d",
                 2623,
                 
                 P
                 , 
                 
                 366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000000; B = 6'b010110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000000; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2624,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b011011; B = 6'b101011; // Expected: {'P': 1161}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b011011; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2625,
                 
                 P
                 , 
                 
                 1161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b011011; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2626,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b011110; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b011110; | Outputs: P=%b | Expected: P=%d",
                 2627,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b010010; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2628,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010100; B = 6'b010010; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010100; B = 6'b010010; | Outputs: P=%b | Expected: P=%d",
                 2629,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111001; B = 6'b000011; // Expected: {'P': 171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111001; B = 6'b000011; | Outputs: P=%b | Expected: P=%d",
                 2630,
                 
                 P
                 , 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110110; B = 6'b110000; // Expected: {'P': 2592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110110; B = 6'b110000; | Outputs: P=%b | Expected: P=%d",
                 2631,
                 
                 P
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b010101; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b010101; | Outputs: P=%b | Expected: P=%d",
                 2632,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b010011; // Expected: {'P': 342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b010011; | Outputs: P=%b | Expected: P=%d",
                 2633,
                 
                 P
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111100; B = 6'b010100; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111100; B = 6'b010100; | Outputs: P=%b | Expected: P=%d",
                 2634,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b110101; B = 6'b011111; // Expected: {'P': 1643}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b110101; B = 6'b011111; | Outputs: P=%b | Expected: P=%d",
                 2635,
                 
                 P
                 , 
                 
                 1643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b000100; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b000100; | Outputs: P=%b | Expected: P=%d",
                 2636,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b000001; // Expected: {'P': 61}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b000001; | Outputs: P=%b | Expected: P=%d",
                 2637,
                 
                 P
                 , 
                 
                 61
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000110; B = 6'b100111; // Expected: {'P': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000110; B = 6'b100111; | Outputs: P=%b | Expected: P=%d",
                 2638,
                 
                 P
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101011; B = 6'b011010; // Expected: {'P': 1118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101011; B = 6'b011010; | Outputs: P=%b | Expected: P=%d",
                 2639,
                 
                 P
                 , 
                 
                 1118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b001010; B = 6'b100100; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b001010; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2640,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101010; B = 6'b001011; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101010; B = 6'b001011; | Outputs: P=%b | Expected: P=%d",
                 2641,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111011; B = 6'b100101; // Expected: {'P': 2183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111011; B = 6'b100101; | Outputs: P=%b | Expected: P=%d",
                 2642,
                 
                 P
                 , 
                 
                 2183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111000; B = 6'b110100; // Expected: {'P': 2912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111000; B = 6'b110100; | Outputs: P=%b | Expected: P=%d",
                 2643,
                 
                 P
                 , 
                 
                 2912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b011011; // Expected: {'P': 1026}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b011011; | Outputs: P=%b | Expected: P=%d",
                 2644,
                 
                 P
                 , 
                 
                 1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010110; B = 6'b010111; // Expected: {'P': 506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010110; B = 6'b010111; | Outputs: P=%b | Expected: P=%d",
                 2645,
                 
                 P
                 , 
                 
                 506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100010; B = 6'b010110; // Expected: {'P': 748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100010; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2646,
                 
                 P
                 , 
                 
                 748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101101; B = 6'b101011; // Expected: {'P': 1935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101101; B = 6'b101011; | Outputs: P=%b | Expected: P=%d",
                 2647,
                 
                 P
                 , 
                 
                 1935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b111101; B = 6'b100010; // Expected: {'P': 2074}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b111101; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 2648,
                 
                 P
                 , 
                 
                 2074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b100100; // Expected: {'P': 1584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b100100; | Outputs: P=%b | Expected: P=%d",
                 2649,
                 
                 P
                 , 
                 
                 1584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101100; B = 6'b100010; // Expected: {'P': 1496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101100; B = 6'b100010; | Outputs: P=%b | Expected: P=%d",
                 2650,
                 
                 P
                 , 
                 
                 1496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010001; B = 6'b111011; // Expected: {'P': 1003}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010001; B = 6'b111011; | Outputs: P=%b | Expected: P=%d",
                 2651,
                 
                 P
                 , 
                 
                 1003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000010; B = 6'b010110; // Expected: {'P': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000010; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2652,
                 
                 P
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100101; B = 6'b100000; // Expected: {'P': 1184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100101; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2653,
                 
                 P
                 , 
                 
                 1184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100001; B = 6'b010110; // Expected: {'P': 726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100001; B = 6'b010110; | Outputs: P=%b | Expected: P=%d",
                 2654,
                 
                 P
                 , 
                 
                 726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b000011; B = 6'b111110; // Expected: {'P': 186}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b000011; B = 6'b111110; | Outputs: P=%b | Expected: P=%d",
                 2655,
                 
                 P
                 , 
                 
                 186
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b010010; B = 6'b111010; // Expected: {'P': 1044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b010010; B = 6'b111010; | Outputs: P=%b | Expected: P=%d",
                 2656,
                 
                 P
                 , 
                 
                 1044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b101110; B = 6'b100000; // Expected: {'P': 1472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b101110; B = 6'b100000; | Outputs: P=%b | Expected: P=%d",
                 2657,
                 
                 P
                 , 
                 
                 1472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100000; B = 6'b110101; // Expected: {'P': 1696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100000; B = 6'b110101; | Outputs: P=%b | Expected: P=%d",
                 2658,
                 
                 P
                 , 
                 
                 1696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 6'b100110; B = 6'b001100; // Expected: {'P': 456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 6'b100110; B = 6'b001100; | Outputs: P=%b | Expected: P=%d",
                 2659,
                 
                 P
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule