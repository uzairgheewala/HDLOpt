
`timescale 1ns / 1ps

module tb_N64_kogge_stone_adder;

    // Parameters
    
    parameter N = 64;
    
     
    // Inputs
    
    reg  [63:0] a;
    
    reg  [63:0] b;
    
    
    // Outputs
    
    wire  [63:0] sum;
    
    wire   cout;
    
    
    // Instantiate the Unit Under Test (UUT)
    kogge_stone_adder  #( N ) uut (
        
        .a(a),
        
        .b(b),
        
        
        .sum(sum),
        
        .cout(cout)
        
    );
    
    initial begin
        // Initialize Inputs
        
        a = 0;
        
        b = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        a = 64'b0000000000000000000000000000000000000000000000001011110110101000; b = 64'b0000000000000000000000000000000000000000000000001110111111110100; // Expected: {'sum': 109980, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001011110110101000; b = 64'b0000000000000000000000000000000000000000000000001110111111110100; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 0,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 109980, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001011101011101100; b = 64'b0000000000000000000000000000000000000000000000000111111101100100; // Expected: {'sum': 80464, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001011101011101100; b = 64'b0000000000000000000000000000000000000000000000000111111101100100; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 1,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 80464, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000000011011100010; b = 64'b0000000000000000000000000000000000000000000000001010010110011101; // Expected: {'sum': 44159, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000000011011100010; b = 64'b0000000000000000000000000000000000000000000000001010010110011101; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 2,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 44159, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001100010010111101; b = 64'b0000000000000000000000000000000000000000000000001110101110000001; // Expected: {'sum': 110654, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001100010010111101; b = 64'b0000000000000000000000000000000000000000000000001110101110000001; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 3,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 110654, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000110100010010010; b = 64'b0000000000000000000000000000000000000000000000000011000010101000; // Expected: {'sum': 39226, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000110100010010010; b = 64'b0000000000000000000000000000000000000000000000000011000010101000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 4,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 39226, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001100010011110010; b = 64'b0000000000000000000000000000000000000000000000001000110101110010; // Expected: {'sum': 86628, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001100010011110010; b = 64'b0000000000000000000000000000000000000000000000001000110101110010; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 5,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 86628, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000010000100101010; b = 64'b0000000000000000000000000000000000000000000000001011000000011100; // Expected: {'sum': 53574, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000010000100101010; b = 64'b0000000000000000000000000000000000000000000000001011000000011100; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 6,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 53574, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001001000011010101; b = 64'b0000000000000000000000000000000000000000000000000101011000000100; // Expected: {'sum': 59097, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001001000011010101; b = 64'b0000000000000000000000000000000000000000000000000101011000000100; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 7,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59097, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000001110111100100; b = 64'b0000000000000000000000000000000000000000000000001110011001100111; // Expected: {'sum': 66635, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000001110111100100; b = 64'b0000000000000000000000000000000000000000000000001110011001100111; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 8,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 66635, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001100110101100110; b = 64'b0000000000000000000000000000000000000000000000000000111011000010; // Expected: {'sum': 56360, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001100110101100110; b = 64'b0000000000000000000000000000000000000000000000000000111011000010; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 9,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 56360, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000000110010111101; b = 64'b0000000000000000000000000000000000000000000000000001110000110111; // Expected: {'sum': 10484, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000000110010111101; b = 64'b0000000000000000000000000000000000000000000000000001110000110111; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 10,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 10484, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000111100001000100; b = 64'b0000000000000000000000000000000000000000000000000001110001001111; // Expected: {'sum': 38035, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000111100001000100; b = 64'b0000000000000000000000000000000000000000000000000001110001001111; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 11,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 38035, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000100001011101101; b = 64'b0000000000000000000000000000000000000000000000000101111100100011; // Expected: {'sum': 41488, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000100001011101101; b = 64'b0000000000000000000000000000000000000000000000000101111100100011; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 12,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 41488, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000011001111100100; b = 64'b0000000000000000000000000000000000000000000000001000011001000000; // Expected: {'sum': 47652, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000011001111100100; b = 64'b0000000000000000000000000000000000000000000000001000011001000000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 13,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 47652, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000010000110001011; b = 64'b0000000000000000000000000000000000000000000000001010001011000111; // Expected: {'sum': 50258, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000010000110001011; b = 64'b0000000000000000000000000000000000000000000000001010001011000111; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 14,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50258, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001100100101100111; b = 64'b0000000000000000000000000000000000000000000000001001101011100110; // Expected: {'sum': 91213, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001100100101100111; b = 64'b0000000000000000000000000000000000000000000000001001101011100110; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 15,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 91213, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001000011011010011; b = 64'b0000000000000000000000000000000000000000000000000000000110000010; // Expected: {'sum': 34901, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001000011011010011; b = 64'b0000000000000000000000000000000000000000000000000000000110000010; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 16,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 34901, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001101101110010010; b = 64'b0000000000000000000000000000000000000000000000001011011101101110; // Expected: {'sum': 103168, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001101101110010010; b = 64'b0000000000000000000000000000000000000000000000001011011101101110; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 17,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 103168, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000001110011010010; b = 64'b0000000000000000000000000000000000000000000000000110001100101100; // Expected: {'sum': 32766, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000001110011010010; b = 64'b0000000000000000000000000000000000000000000000000110001100101100; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 18,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 32766, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001000100110100110; b = 64'b0000000000000000000000000000000000000000000000001000011100100010; // Expected: {'sum': 69832, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001000100110100110; b = 64'b0000000000000000000000000000000000000000000000001000011100100010; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 19,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69832, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001101000111101000; b = 64'b0000000000000000000000000000000000000000000000000111100001101010; // Expected: {'sum': 84562, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001101000111101000; b = 64'b0000000000000000000000000000000000000000000000000111100001101010; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 20,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 84562, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000000000100111011; b = 64'b0000000000000000000000000000000000000000000000001110010110001000; // Expected: {'sum': 59075, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000000000100111011; b = 64'b0000000000000000000000000000000000000000000000001110010110001000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 21,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 59075, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001000110100000101; b = 64'b0000000000000000000000000000000000000000000000000010100100011101; // Expected: {'sum': 46626, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001000110100000101; b = 64'b0000000000000000000000000000000000000000000000000010100100011101; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 22,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 46626, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000110010010111101; b = 64'b0000000000000000000000000000000000000000000000000101100111100001; // Expected: {'sum': 48798, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000110010010111101; b = 64'b0000000000000000000000000000000000000000000000000101100111100001; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 23,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 48798, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000101111100110111; b = 64'b0000000000000000000000000000000000000000000000000111011010111011; // Expected: {'sum': 54770, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000101111100110111; b = 64'b0000000000000000000000000000000000000000000000000111011010111011; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 24,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 54770, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000111101010001111; b = 64'b0000000000000000000000000000000000000000000000001001010101010110; // Expected: {'sum': 69605, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000111101010001111; b = 64'b0000000000000000000000000000000000000000000000001001010101010110; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 25,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 69605, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001110010111011011; b = 64'b0000000000000000000000000000000000000000000000000111010010001110; // Expected: {'sum': 88681, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001110010111011011; b = 64'b0000000000000000000000000000000000000000000000000111010010001110; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 26,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 88681, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001101000010111010; b = 64'b0000000000000000000000000000000000000000000000000110110011101010; // Expected: {'sum': 81316, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001101000010111010; b = 64'b0000000000000000000000000000000000000000000000000110110011101010; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 27,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 81316, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001110110011110100; b = 64'b0000000000000000000000000000000000000000000000000101001101100000; // Expected: {'sum': 82004, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001110110011110100; b = 64'b0000000000000000000000000000000000000000000000000101001101100000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 28,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 82004, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000111011001100011; b = 64'b0000000000000000000000000000000000000000000000000110000010100000; // Expected: {'sum': 55043, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000111011001100011; b = 64'b0000000000000000000000000000000000000000000000000110000010100000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 29,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 55043, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001100100111100000; b = 64'b0000000000000000000000000000000000000000000000001001100001000000; // Expected: {'sum': 90656, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001100100111100000; b = 64'b0000000000000000000000000000000000000000000000001001100001000000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 30,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 90656, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000001010100010100100; b = 64'b0000000000000000000000000000000000000000000000000111010100010000; // Expected: {'sum': 73140, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000001010100010100100; b = 64'b0000000000000000000000000000000000000000000000000111010100010000; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 31,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 73140, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        a = 64'b0000000000000000000000000000000000000000000000000111101101010011; b = 64'b0000000000000000000000000000000000000000000000000100100101100101; // Expected: {'sum': 50360, 'cout': 0}
        #10;
        $display("Test %0d: Inputs: a = 64'b0000000000000000000000000000000000000000000000000111101101010011; b = 64'b0000000000000000000000000000000000000000000000000100100101100101; | Outputs: sum=%b, cout=%b | Expected: sum=%d, cout=%d",
                 32,
                 
                 sum, 
                 
                 cout
                 , 
                 
                 50360, 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule